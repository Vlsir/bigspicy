** Translated using xdm 2.6.0 on Nov_14_2022_16_05_33_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 2
.PARAM 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__TOXE_MULT=1.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__RBPB_MULT=1.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__OVERLAP_MULT=0.89805 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__AJUNCTION_MULT=9.9505e-1 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__PJUNCTION_MULT=1.0144 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__LINT_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__WINT_DIFF=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__RSHG_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__DLC_DIFF=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__XGW_DIFF=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VTH0_DIFF_0=-0.015262 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VSAT_DIFF_0=-3503.4 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__K2_DIFF_0=0.0013127 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__U0_DIFF_0=-0.0029685 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VTH0_DIFF_1=-0.0025365 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VSAT_DIFF_1=323.35 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__K2_DIFF_1=-0.00053421 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__U0_DIFF_1=-0.0010115 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VSAT_DIFF_0=-3946.4 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VTH0_DIFF_0=-0.024526 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__K2_DIFF_0=0.0010173 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__U0_DIFF_0=-0.0031271 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VSAT_DIFF_1=-1841.7 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VTH0_DIFF_1=-0.0099998 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__K2_DIFF_1=-0.00057848 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__U0_DIFF_1=-0.0013993 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VSAT_DIFF_2=-2994.9 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VTH0_DIFF_2=-0.0082165 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__K2_DIFF_2=-0.0015137 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__U0_DIFF_2=-0.003002 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__K2_DIFF_0=0.00059498 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__U0_DIFF_0=-0.0016449 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VTH0_DIFF_0=-0.015075 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VSAT_DIFF_0=1100.9 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__K2_DIFF_1=-0.0068059 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__U0_DIFF_1=-0.002939 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VTH0_DIFF_1=-0.012671 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VSAT_DIFF_1=-3862.9 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__K2_DIFF_2=-0.0017173 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__U0_DIFF_2=-0.0041054 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VTH0_DIFF_2=-0.022123 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VSAT_DIFF_2=-5556.8
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
*





* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 002, W = 7.09, L = 0.5
* --------------------------------------------
*















* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 000, W = 3.01, L = 0.5
* ---------------------------------------------
*















* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 001, W = 5.05, L = 0.5
* ---------------------------------------------
*















* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 002, W = 7.09, L = 0.5
* ---------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice















