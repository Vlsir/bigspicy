** Translated using xdm 2.6.0 on Nov_14_2022_16_05_26_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__cap_var_hvt c0 c1 b 
+ PARAMS: W=5 L=0.5 VM=1 WC='w*1' LC='l*1'
* Corner Parameters
*.param cnwvc2_tox=41.7642
*.param cnwvc2_cdepmult=1
*.param cnwvc2_cintmult=1
*.param cnwvc2_vt1=0.2
*.param cnwvc2_vt2=0.33
*.param cnwvc2_vtr=0.14
*.param cnwvc2_dwc=0.0
*.param cnwvc2_dlc=0.0
*.param cnwvc2_dld=0.0
* Geometry Parameters
.PARAM 
+ CNWVC_LDIFF=0.15 WD='wc+2*cnwvc2_dwc' LD='lc+2*cnwvc2_dlc' LDD='0.015+2*cnwvc2_dld' 
+ DWR=0.00 DWP=0.0 DLR=0.03 WL='(wd-2*dwr)/(ld-2*dlr)' WLWDIFF='((0.5*(ld-2*dlr))+cnwvc_ldiff)/(2*(wd-2*dwr))' 
+ SKY130_FD_PR__CAP_VAR_HVT__CMIN_SLOPE_L=2.4e-16 SKY130_FD_PR__CAP_VAR_HVT__CMIN_SLOPE_W=1.0e-16 
+ SKY130_FD_PR__CAP_VAR_HVT__CMIN_SLOPE_WL=4.0e-16 SKY130_FD_PR__CAP_VAR_HVT__CMAX_SLOPE_L=3.0e-16 
+ SKY130_FD_PR__CAP_VAR_HVT__CMAX_SLOPE_W=7.0e-16 SKY130_FD_PR__CAP_VAR_HVT__CMAX_SLOPE_WL=1.0e-15
* Mismatch Parameters




* Capacitance Model Parameters






.PARAM CNWVC_SLOPE1=0.15
.PARAM CNWVC_SLOPE2=0.35
.PARAM 
+ CM0='5.828e-16*cnwvc2_cintmult' CM1='4.596e-16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*sky130_fd_pr__cap_var_hvt__cmin_slope_l/sqrt(2*ld*vm)' 
+ CM2='1.614e-16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*sky130_fd_pr__cap_var_hvt__cmin_slope_w/sqrt(2*wd*vm)' 
+ CM3='1.541e-15*cnwvc2_cdepmult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*sky130_fd_pr__cap_var_hvt__cmin_slope_wl*cnwvc2_cdepmult/sqrt(2*ld*wd*vm)' 
+ CX0=6.778e-16 CX1='6.461e-16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*sky130_fd_pr__cap_var_hvt__cmax_slope_l/sqrt(2*ld*vm)' 
+ CX2='1.517e-16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*sky130_fd_pr__cap_var_hvt__cmax_slope_w/sqrt(2*wd*vm)' 
+ CX3='8.854e-14*3.9/cnwvc2_tox+MC_MM_SWITCH*AGAUSS(0,1.0,1)*sky130_fd_pr__cap_var_hvt__cmax_slope_wl/sqrt(2*ld*wd*vm)' 
+ SKY130_FD_PR__CAP_VAR_HVT__VGS_MIN_1='-2.071' SKY130_FD_PR__CAP_VAR_HVT__VGS_MAX_1='-1*-2.071' 
+ SKY130_FD_PR__CAP_VAR_HVT__TMAX_VGS_1='100.001n' SKY130_FD_PR__CAP_VAR_HVT__VGS_MIN_2='-2.161' 
+ SKY130_FD_PR__CAP_VAR_HVT__VGS_MAX_2='-1*-2.161' SKY130_FD_PR__CAP_VAR_HVT__TMAX_VGS_2='20.001n' 
+ SKY130_FD_PR__CAP_VAR_HVT__VGS_MIN='-2.301' SKY130_FD_PR__CAP_VAR_HVT__VGS_MAX='-1*-2.301'
* .SETSOA LABEL="MODEL_OOB_VG_1: sky130_fd_pr__cap_var_hvt Vg for Varactor" E v(c0, c1) =(sky130_fd_pr__cap_var_hvt__vgs_min_1, sky130_fd_pr__cap_var_hvt__vgs_max_1, sky130_fd_pr__cap_var_hvt__tmax_vgs_1 )






* .SETSOA LABEL="MODEL_OOB_VG_2: sky130_fd_pr__cap_var_hvt Vg for Varactor" E v(c0, c1) =(sky130_fd_pr__cap_var_hvt__vgs_min_2, sky130_fd_pr__cap_var_hvt__vgs_max_2, sky130_fd_pr__cap_var_hvt__tmax_vgs_2 )
* .SETSOA LABEL="MODEL_OOB_VG: sky130_fd_pr__cap_var_hvt Vg for Varactor" E v(c0, c1) =(sky130_fd_pr__cap_var_hvt__vgs_min, sky130_fd_pr__cap_var_hvt__vgs_max )
.PARAM 
+ TREF=30.0 CMIN='cm0+cm1*ld+cm2*wd+cm3*wd*(ld-ldd)+cx3*wd*ldd' CMAX='cx0+cx1*ld+cx2*wd+cx3*wd*ld' 
+ SLOPE_0=1.808e-17 SLOPE_0_TC1=7.2181e-20 SLOPE_0_TC2=-1.9745e-21 CMIN_SLOPE_0='slope_0+(temp-tref)*slope_0_tc1+(temp-tref)*(temp-tref)*slope_0_tc2' 
+ SLOPE_W=-3.169e-17 SLOPE_W_TC1=-1.4465e-19 SLOPE_W_TC2=3.5187e-21 CMIN_SLOPE_W='slope_w+(temp-tref)*slope_w_tc1+(temp-tref)*(temp-tref)*slope_w_tc2' 
+ SLOPE_L=-7.435e-17 SLOPE_L_TC1=-4.4474e-19 SLOPE_L_TC2=7.3824e-21 CMIN_SLOPE_L='slope_l+(temp-tref)*slope_l_tc1+(temp-tref)*(temp-tref)*slope_l_tc2' 
+ SLOPE_WL=2.509e-16 SLOPE_WL_TC1=-1.0793e-18 SLOPE_WL_TC2=-2.2625e-20 CMIN_SLOPE_WL='slope_wl+(temp-tref)*slope_wl_tc1+(temp-tref)*(temp-tref)*slope_wl_tc2' 
+ CMIN_SLOPE='cmin_slope_0+cmin_slope_w*wd+cmin_slope_l*ld+cmin_slope_wl*wd*ld'
Cg c0 p2














C3 c0 b C='0.15e-15'
C4 c1 b C='0.15e-15'
* Resistance Model Parameters
.PARAM CON_SP=0.17
.PARAM CNWVC_K=12
.PARAM CNWVC_N1=0.2
.PARAM CNWVC_N2=0.35
.PARAM APOLY=1.1
.PARAM APOLYC=1.1
.PARAM ACON=1
.PARAM ANWELL=1
.PARAM BNWELL=0.5
.PARAM CNWELL=0.3
.PARAM N_POCON='max((lc-0.14)/(2*con_sp),1)'
.PARAM N_CON='(wc-2*0.06+con_sp)/(2*con_sp)'
.PARAM RG_TC1=9.611e-4
.PARAM RG_TC2=5.523e-6
.PARAM RG_TCMULT='1+(temp-tref)*rg_tc1+(temp-tref)*(temp-tref)*rg_tc2'
.PARAM 
+ CNWVC_A='apoly*rp1*wl/cnwvc_k+apolyc*rcp1/n_pocon+acon*rcn/n_con+anwell*rnw*wlwdiff'
.PARAM CNWVC_B1='bnwell*rnw*cnwvc_ldiff/(2*(wd-2*dwr))'
.PARAM CNWVC_C='cnwell*rnw*cnwvc_ldiff/(2*(wd-2*dwp))'
Rg p2 c1 
+ R='(cnwvc_a+cnwvc_b1*(0.5*tanh((v(c0)-v(p2)-cnwvc2_vtr)/cnwvc_n1)+0.5)+20*cnwvc_c*(0.5*tanh((v(c0)-v(p2)-cnwvc2_vtr)/cnwvc_n1)+0.5)*exp(-abs((v(c0)-v(p2)-cnwvc2_vtr)/cnwvc_n2)))/vm*rg_tcmult'
.ENDS sky130_fd_pr__cap_var_hvt
