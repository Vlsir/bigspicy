** Translated using xdm 2.6.0 on Nov_14_2022_16_05_20_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__RF_PFET_01V8_B__TOXE_MULT=0.9635 SKY130_FD_PR__RF_PFET_01V8_B__RBPB_MULT=0.8 
+ SKY130_FD_PR__RF_PFET_01V8_B__OVERLAP_MULT=0.88516 SKY130_FD_PR__RF_PFET_01V8_B__AJUNCTION_MULT=0.93001 
+ SKY130_FD_PR__RF_PFET_01V8_B__PJUNCTION_MULT=0.93439 SKY130_FD_PR__RF_PFET_01V8_B__LINT_DIFF=1.21275e-8 
+ SKY130_FD_PR__RF_PFET_01V8_B__WINT_DIFF=-2.252e-8 SKY130_FD_PR__RF_PFET_01V8_B__RSHG_DIFF=-7.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__DLC_DIFF=1.21275e-8 SKY130_FD_PR__RF_PFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__XGW_DIFF=-4.504e-8 SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT=0.8875 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT=0.839 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT=0.839 
+ SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT_2=0.8875 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT_2=0.86 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT_2=0.86 SKY130_FD_PR__RF_PFET_01V8__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RS_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_0=-0.0096187 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_0=-9.1722e-5 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_0=-0.057483 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_0=-11003.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_1=-0.012861 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_1=1.6284e-5 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_1=-0.054689 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_1=-6396.5 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_2=-0.029824 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_2=0.00016037 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_2=-0.02191 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_2=5271.4 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_3=-0.013607 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_3=3.7455e-6 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_3=-0.077102 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_3=-10440.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_4=-0.0077158 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_4=-0.00015599 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_4=-0.04551 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_4=-2665.7 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_5=-0.018523 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_5=2.6323e-5 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_5=-0.017911 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_5=11962.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_6=-0.013977 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_6=-0.00029174 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_6=-0.081869 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_6=-8538.5 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_7=-3.0985e-5 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_7=-8661.9 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_7=-0.0068507 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_7=-0.050877 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_8=-0.024781 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_8=-3.1187e-5 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_8=3310.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_8=-0.020378 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_0=-0.007218 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_0=-0.00024908 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_0=-0.045584 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_0=-10840.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_1=-0.011746 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_1=-5.8756e-5 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_1=-0.040864 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_1=-2721.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_2=0.00011377 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_2=-0.014596 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_2=11806.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_2=-0.030918 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_3=-0.011489 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_3=-0.00010472 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_3=-0.075251 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_3=-6951.2 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_4=-0.00033553 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_4=-0.032126 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_4=-3166.2 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_4=-0.0039733 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_5=-0.0099782 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_5=-7.0926e-5 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_5=7638.8 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_5=-0.018384 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_6=-0.076598 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_6=-0.00010558 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_6=-8165.2 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_6=-0.012381 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_7=-0.0043219 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_7=-0.046792 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_7=-0.00030508 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_7=-6293.3 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_8=-0.018996 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_8=-0.012116 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_8=-0.00013862 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_8=17138.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_8=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_pfet_01v8_b.pm3.spice














