** Translated using xdm 2.6.0 on Nov_14_2022_16_05_20_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__TOXE_MULT=0.9635 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RBPB_MULT=0.8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__OVERLAP_MULT=8.8119e-1 SKY130_FD_PR__RF_NFET_01V8_LVT_B__AJUNCTION_MULT=8.7784e-1 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__PJUNCTION_MULT=7.8244e-1 SKY130_FD_PR__RF_NFET_01V8_LVT_B__LINT_DIFF=1.21275e-8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__WINT_DIFF=-2.252e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RSHG_DIFF=-7.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__DLC_DIFF=7.7131e-9 SKY130_FD_PR__RF_NFET_01V8_LVT_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__XGW_DIFF=-4.504e-8 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT_P42=0.8875 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT_P42=0.755 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT_P42=0.755 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT=0.8875 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT=0.825 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT=0.825 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RS_MULT=1.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_0=-0.043187 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_0=0.0031893 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_0=-20156.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_0=-0.0091082 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_1=-0.00023031 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_1=-0.039728 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_1=0.0032163 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_1=-16799.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_2=-0.0031116 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_2=-0.032085 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_2=0.003301 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_2=-12923.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_3=0.0056278 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_3=-0.051298 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_3=-0.001719 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_3=-25716.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_4=0.0040629 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_4=-0.050969 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_4=-0.001606 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_4=-16982.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_5=0.0028518 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_5=-0.021748 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_5=0.001153 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_5=-11783.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_6=-0.0053048 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_6=-0.045076 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_6=-0.0074793 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_6=-20834.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_7=0.0027467 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_7=-0.042761 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_7=-0.0034925 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_7=-14000.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_8=0.0026278 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_8=-0.018088 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_8=0.00072051 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_8=-10215.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_0=-0.0093685 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_0=-0.046477 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_0=-0.003305 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_0=-16286.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_1=-0.0011171 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_1=-0.047694 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_1=-0.00091767 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_1=-16903.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_2=0.0014264 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_2=-0.037401 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_2=0.00086418 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_2=-7635.6 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_3=0.004034 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_3=-0.049369 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_3=-0.0026239 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_3=-26112.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_4=-0.0064811 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_4=-15470.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_4=0.002107 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_4=-0.046682 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_5=-0.033495 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_5=-0.002231 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_5=-2766.3 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_5=0.0013838 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_6=-0.0022088 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_6=-0.049429 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_6=-0.0050469 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_6=-24301.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_7=-0.00079282 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_7=-0.042712 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_7=-0.0075496 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_7=-16463.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_8=0.00082322 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_8=-0.0041644 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_8=-543.48 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_8=-0.034543 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_8=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice















