** Translated using xdm 2.6.0 on Nov_14_2022_16_05_11_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
