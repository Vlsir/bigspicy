** Translated using xdm 2.6.0 on Nov_14_2022_16_05_30_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65 l = 0.15 m = 2 ad = 0.231 pd = 1.93 as = 0.462 ps = 3.86 nrd = 240.00 nrs = 120.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65 l = 0.15 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 120.0 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65 l = 0.15 m = 4 ad = 0.231 pd = 1.93 as = 0.347 ps = 2.90 nrd = 240.00 nrs = 160.00 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65 l = 0.15 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 120.00 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65 l = 0.18 m = 2 ad = 0.231 pd = 1.93 as = 0.462 ps = 3.86 nrd = 240.00 nrs = 120.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65 l = 0.18 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 120.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65 l = 0.18 m = 4 ad = 0.231 pd = 1.93 as = 0.347 ps = 2.90 nrd = 240.00 nrs = 160.00 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65 l = 0.18 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 120.00 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65 l = 0.25 m = 2 ad = 0.231 pd = 1.93 as = 0.462 ps = 3.86 nrd = 240.00 nrs = 120.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65 l = 0.25 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 120.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65 l = 0.25 m = 4 ad = 0.231 pd = 1.93 as = 0.347 ps = 2.90 nrd = 240.00 nrs = 160.00 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65 l = 0.25 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 120.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.15 m = 2 ad = 0.421 pd = 3.29 as = 0.843 ps = 6.58 nrd = 133.33 nrs = 66.67 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.15 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 66.67 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.15 m = 4 ad = 0.421 pd = 3.29 as = 0.632 ps = 4.94 nrd = 133.33 nrs = 88.89 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.15 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 66.67 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.18 m = 2 ad = 0.421 pd = 3.29 as = 0.843 ps = 6.58 nrd = 133.33 nrs = 66.67 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.18 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 66.67 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.18 m = 4 ad = 0.421 pd = 3.29 as = 0.632 ps = 4.94 nrd = 133.33 nrs = 88.89 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.18 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 66.67 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.25 m = 2 ad = 0.421 pd = 3.29 as = 0.843 ps = 6.58 nrd = 133.33 nrs = 66.67 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.25 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 66.67 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.25 m = 4 ad = 0.421 pd = 3.29 as = 0.632 ps = 4.94 nrd = 133.33 nrs = 88.89 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.25 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 66.67 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.15 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 80.00 nrs = 40.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.15 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 40.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.15 m = 4 ad = 0.707 pd = 5.33 as = 1.061 ps = 8.00 nrd = 80.00 nrs = 53.33 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.15 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 40.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.18 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 80.00 nrs = 40.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.18 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 40.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.18 m = 4 ad = 0.707 pd = 5.33 as = 1.061 ps = 8.00 nrd = 80.00 nrs = 53.33 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.18 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 40.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.25 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 80.00 nrs = 40.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.25 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 40.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25
.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.25 m = 4 ad = 0.707 pd = 5.33 as = 1.061 ps = 8.00 nrd = 80.00 nrs = 53.33 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.25 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 40.00 nrs = 0.00 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25
.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 d g s b
* .param  mult = 1.0  rg_sub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult)}   rg_dist_tnom = {(150.129*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15 w = {(2)*(1.68)} ad = {(2)*(0.2352)} as = {(2)*(0.445)} pd = {(2)*(1.96)} ps = {(2)*(3.89)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(0.41f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(0.74f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.119f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_sub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(154*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(76*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 d g s b
* .param  mult = 1.0  rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2)}   rg_dist_tnom = {(366.81*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15 w = {(2)*(5.00)} ad = {(2)*(0.7)} as = {(2)*(1.325)} pd = {(2)*(5.28)} ps = {(2)*(10.53)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(1.22f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(1.665f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.285f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(50*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(24*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15 d g s b
* .param  mult = 1.0  rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2)}   rg_dist_tnom = {(37.53*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15 w = {(2)*(0.84)} ad = {(2)*(0.1176)} as = {(2)*(0.223)} pd = {(2)*(1.12)} ps = {(2)*(2.21)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(0.17f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(0.459f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.257f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(306*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(152.5*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15 d g s b
* .param  mult = 1.0  rg_stub_tnom = {(63.5*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult)}   rg_dist_tnom = {(75.061*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15 w = {(4)*(1.68)} ad = {(4)*(0.2352)} as = {(4)*(0.34)} pd = {(4)*(1.96)} ps = {(4)*(2.925)} nrd = {(0)/(4)} nrs = {(0)/(4)} nf = 4 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(0.82f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(0.984f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.354f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(78*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(50.6*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 d g s b
* .param  mult = 1.0  rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult)}   rg_dist_tnom = {(183.0*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15 w = {(2)*(3.00)} ad = {(2)*(0.42)} as = {(2)*(0.795)} pd = {(2)*(3.28)} ps = {(2)*(6.53)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3  c = {(0.7f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1  c = {(1.056f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3  c = {(0.232f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g  r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d  r = {(78*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s  r = {(38.5*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15
