** Translated using xdm 2.6.0 on Nov_14_2022_16_05_32_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_B__TOXE_MULT=0.948 SKY130_FD_PR__RF_NFET_01V8_B__RBPB_MULT=0.8 
+ SKY130_FD_PR__RF_NFET_01V8_B__OVERLAP_MULT=0.94816 SKY130_FD_PR__RF_NFET_01V8_B__AJUNCTION_MULT=0.7739 
+ SKY130_FD_PR__RF_NFET_01V8_B__PJUNCTION_MULT=0.79336 SKY130_FD_PR__RF_NFET_01V8_B__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__RF_NFET_01V8_B__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__RF_NFET_01V8_B__RSHG_DIFF=-7.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__DLC_DIFF=12.773e-9 SKY130_FD_PR__RF_NFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__XGW_DIFF=-6.4250e-8 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_0=-0.075991 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_0=-22417.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_0=0.010085 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_0=0.00074749 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_1=-0.039487 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_1=-19233.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_1=0.020683 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_1=0.0011292 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_2=-0.043022 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_2=-16781.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_2=0.038033 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_2=0.0006468 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_3=-0.035105 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_3=-28463.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_3=0.010626 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_3=-0.0036794 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_4=-0.05182 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_4=-25171.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_4=0.030375 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_4=-0.0033229 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_5=-0.032322 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_5=-20257.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_5=0.042979 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_5=0.0011015 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_6=-0.0033456 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_6=-0.041439 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_6=-28660.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_6=0.0064952 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_7=0.02645 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_7=-0.0036669 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_7=-0.045761 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_7=-23039.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_8=0.04175 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_8=-0.0010573 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_8=-0.032973 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_8=-16043.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_0=0.0091842 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_0=-0.00070926 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_0=-0.051501 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_0=-31984.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_1=0.028977 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_1=-0.0013648 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_1=-0.058125 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_1=-23564.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_2=0.042169 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_2=-0.00035031 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_2=-0.046633 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_2=-19030.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_3=-30928.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_3=0.013856 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_3=-0.0048131 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_3=-0.046817 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_4=-24921.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_4=0.034977 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_4=-0.0071423 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_4=-0.061148 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_5=-8528.2 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_5=0.045401 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_5=-0.0043436 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_5=-0.04118 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_6=-29958.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_6=0.009601 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_6=-0.0033405 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_6=-0.04502 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_7=-0.0060347 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_7=-26996.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_7=0.031931 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_7=-0.060436 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_8=-0.0389 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_8=-0.0030982 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_8=-11896.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_8=0.044114
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*





* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_b.pm3.spice














