** Translated using xdm 2.6.0 on Nov_14_2022_16_05_20_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_01V8_LVT__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__nfet_01v8_lvt d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__nfet_01v8_lvt d g s b sky130_fd_pr__nfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__nfet_01v8_lvt__model.0 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.417702+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47213   k2 = -0.0340947   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 161140.0   ua = -1.3015598e-9   ub = 2.68715e-18   uc = 7.0152e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0321123   a0 = 1.95580301   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.554525   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11559919+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.0383479+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0047977   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.4345657e-5   alpha1 = 0.0   beta0 = 17.822982   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25364   kt2 = -0.034423   at = 333080.0   ute = -1.0777   ua1 = 2.6823e-9   ub1 = -2.4433e-18   uc1 = -1.9223e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.1 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.082993200e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = 7.476724334e-08 wvth0 = 6.575331717e-08 pvth0 = -5.228503233e-13   k1 = 5.484178983e-01 lk1 = -6.066180995e-07 wk1 = -5.334843243e-07 pk1 = 4.242104634e-12   k2 = -6.014295857e-02 lk2 = 2.071278074e-07 wk2 = 1.821565141e-07 pk2 = -1.448453042e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.424062713e+04 lvsat = 6.909973088e-01 wvsat = 6.076907905e-01 pvsat = -4.832171820e-6   ua = -1.339578462e-09 lua = 3.023128007e-16 wua = 2.658660208e-16 pua = -2.114085508e-21   ub = 2.692004298e-18 lub = -3.859989856e-26 wub = -3.394630134e-26 pub = 2.699306346e-31   uc = 6.984502141e-11 luc = 2.441000150e-18 wuc = 2.146713586e-18 puc = -1.707001169e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.166786085e-02 lu0 = 3.534044542e-09 wu0 = 3.107980732e-09 pu0 = -2.471371484e-14   a0 = 1.993636486e+00 la0 = -3.008402610e-07 wa0 = -2.645710102e-07 pa0 = 2.103787979e-12   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.343483274e-01 lags = 1.604387469e-07 wags = 1.410962788e-07 pags = -1.121954574e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.120894156e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.790865576e-08 wvoff = -2.454399296e-08 pvoff = 1.951663461e-13   nfactor = {1.107586083e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.505609111e-07 wnfactor = -4.841853811e-07 pnfactor = 3.850094474e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 3.397379306e-01 lpclm = -1.111153404e-06 wpclm = -9.771929379e-07 ppclm = 7.770340199e-12   pdiblc1 = 0.39   pdiblc2 = 2.897088242e-03 lpdiblc2 = 1.511308501e-08 wpdiblc2 = 1.329105404e-08 ppdiblc2 = -1.056864080e-13   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.380464198e-04 lalpha0 = -4.270120873e-10 walpha0 = -3.755315825e-10 palpha0 = 2.986112607e-15   alpha1 = 0.0   beta0 = 1.812212786e+01 lbeta0 = -2.378716637e-06 wbeta0 = -2.091938963e-06 pbeta0 = 1.663446059e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.532257382e-01 lkt1 = -3.294083247e-09 wkt1 = -2.896949130e-09 pkt1 = 2.303565591e-14   kt2 = -3.413939002e-02 lkt2 = -2.255180069e-09 wkt2 = -1.983295943e-09 pkt2 = 1.577056443e-14   at = 6.145496287e+05 lat = -2.238160639e+00 wat = -1.968328372e+00 pat = 1.565154687e-5   ute = -9.510846077e-01 lute = -1.006806982e-06 wute = -8.854265032e-07 pute = 7.040641498e-12   ua1 = 2.424183051e-09 lua1 = 2.052467254e-15 wua1 = 1.805022150e-15 pua1 = -1.435298560e-20   ub1 = -1.561878418e-18 lub1 = -7.008795585e-24 wub1 = -6.163816379e-24 pub1 = 4.901278788e-29   uc1 = -1.098556403e-11 luc1 = -6.550157841e-17 wuc1 = -5.760471923e-17 puc1 = 4.580551579e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.2 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.237652312e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.365067941e-08 wvth0 = -1.315066343e-07 pvth0 = 2.566608407e-13   k1 = 3.602860781e-01 lk1 = 1.368214739e-07 wk1 = 1.066968649e-06 pk1 = -2.082397377e-12   k2 = 3.470276840e-03 lk2 = -4.425229689e-08 wk2 = -3.643130282e-07 pk2 = 7.110279155e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.477945333e+05 lvsat = -7.851737944e-01 wvsat = -1.215381581e+00 pvsat = 2.372054155e-6   ua = -1.299861368e-09 lua = 1.453629628e-16 wua = -5.317320415e-16 pua = 1.037778767e-21   ub = 2.635099381e-18 lub = 1.862709796e-25 wub = 6.789260268e-26 pub = -1.325056532e-31   uc = 6.804041512e-11 luc = 9.572253787e-18 wuc = -4.293427172e-18 puc = 8.379460344e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.092629231e-02 lu0 = 6.464497264e-09 wu0 = -6.215961463e-09 pu0 = 1.213166091e-14   a0 = 1.840206672e+00 la0 = 3.054675683e-07 wa0 = 5.291420204e-07 pa0 = -1.032723836e-12   keta = 1.800731392e-01 lketa = -7.115941237e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.616272718e-01 lags = 3.701061042e-06 wags = -2.821925575e-07 pags = 5.507538035e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.223285511e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.255328484e-08 wvoff = 4.908798591e-08 pvoff = -9.580477667e-14   nfactor = {6.413298149e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.291941651e-06 wnfactor = 9.683707622e-07 pnfactor = -1.889964375e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378214013e-01 letab = 2.680094922e-7   dsub = 8.303355979e-01 ldsub = -1.068283831e-6   voffl = 0.0   minv = 0.0   pclm = -1.088488709e-01 lpclm = 6.615248165e-07 wpclm = 1.954385876e-06 ppclm = -3.814365142e-12   pdiblc1 = 0.39   pdiblc2 = 4.799168520e-03 lpdiblc2 = 7.596643889e-09 wpdiblc2 = -2.658210809e-08 ppdiblc2 = 5.188016745e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.348910763e-05 lalpha0 = 3.693948489e-10 walpha0 = 7.510631650e-10 palpha0 = -1.465846224e-15   alpha1 = 0.0   beta0 = 1.383496396e+01 lbeta0 = 1.456284751e-05 wbeta0 = 4.183877926e-06 pbeta0 = -8.165653629e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.544782820e-01 lkt1 = 1.655587768e-09 wkt1 = 5.793898259e-09 pkt1 = -1.130792226e-14   kt2 = -3.964306084e-02 lkt2 = 1.949364841e-08 wkt2 = 3.966591885e-09 pkt2 = -7.741577549e-15   at = 4.503893511e+04 lat = 1.237192125e-02 wat = 3.936656744e+00 pat = -7.683153284e-6   ute = -1.241640738e+00 lute = 1.413822270e-07 wute = 1.770853006e-06 pute = -3.456164958e-12   ua1 = 2.642495993e-09 lua1 = 1.189761093e-15 wua1 = -3.610044300e-15 pua1 = 7.045705410e-21   ub1 = -2.914608997e-18 lub1 = -1.663216919e-24 wub1 = 1.232763276e-23 pub1 = -2.405977921e-29   uc1 = -2.054783950e-11 luc1 = -2.771438225e-17 wuc1 = 1.152094385e-16 puc1 = -2.248536850e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.3 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.271565445e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.031870199e-9   k1 = 4.290481100e-01 lk1 = 2.618959906e-9   k2 = -1.502755751e-02 lk2 = -8.150166079e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.983806128e+04 lvsat = 5.006671224e-2   ua = -9.566940898e-10 lua = -5.243948992e-16   ub = 2.645230060e-18 lub = 1.664989830e-25   uc = 5.999528613e-11 luc = 2.527389180e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.826786436e-02 lu0 = -7.864012204e-9   a0 = 2.185738384e+00 la0 = -3.689049464e-07 wa0 = -3.388131789e-21   keta = -1.459007000e-01 lketa = -7.539261176e-8   a1 = 0.0   a2 = 0.38689047   ags = 8.887389443e-01 lags = 1.260727550e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.170390794e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.229849331e-9   nfactor = {8.688151836e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.479595944e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.475847500e-05 lcit = -9.287091865e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.889454147e-04 leta0 = -1.735943211e-10   etab = -5.405612409e-04 letab = 7.916317106e-11   dsub = -4.321683872e-02 ldsub = 6.366240922e-7   voffl = 0.0   minv = 0.0   pclm = 2.292529914e-01 lpclm = 1.653102352e-9   pdiblc1 = 0.39   pdiblc2 = 7.056963837e-03 lpdiblc2 = 3.190116056e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.850831459e-04 lalpha0 = -1.157423754e-10   alpha1 = 0.0   beta0 = 2.119942742e+01 lbeta0 = 1.896609901e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.507558811e-01 lkt1 = -5.609403487e-9   kt2 = -4.554545142e-02 lkt2 = 3.101331457e-8   at = 3.150280162e+04 lat = 3.879032530e-2   ute = -1.320519505e+00 lute = 2.953295213e-7   ua1 = 3.273417968e-09 lua1 = -4.160617156e-17   ub1 = -3.904795775e-18 lub1 = 2.693256641e-25   uc1 = 1.013012942e-11 luc1 = -8.758842080e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.4 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.424931113e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.563863729e-9   k1 = 4.336971190e-01 lk1 = -1.805478667e-9   k2 = -1.942855901e-02 lk2 = -3.961754960e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.118593496e+04 lvsat = 4.878394760e-2   ua = -1.239921291e-09 lua = -2.548489882e-16   ub = 2.841201885e-18 lub = -2.000642313e-26   uc = 1.063597291e-10 luc = -1.885091678e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.452171324e-02 lu0 = -4.298818913e-9   a0 = 2.105089053e+00 la0 = -2.921513811e-7   keta = -4.200343856e-01 lketa = 1.854990462e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.012014914e+00 lags = -7.599835742e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.149556753e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.470840543e-10   nfactor = {1.434377196e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.097170550e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 7.647702706e-04 leta0 = -3.409259574e-10   etab = -8.141412672e-04 letab = 3.395279142e-10   dsub = 2.875996857e-01 ldsub = 3.217876600e-7   voffl = 0.0   minv = 0.0   pclm = -2.739760780e-02 lpclm = 2.459061944e-7   pdiblc1 = 0.39   pdiblc2 = 1.030872371e-02 lpdiblc2 = 9.543244381e-11   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.349094263e-05 lalpha0 = 8.275654177e-11 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.870548176e+01 lbeta0 = 2.563136612e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.509857447e-01 lkt1 = -5.390643448e-9   kt2 = -1.928511490e-03 lkt2 = -1.049670907e-8   at = 7.235866273e+04 lat = -9.199343683e-5   ute = -1.005321694e+00 lute = -4.642659429e-9   ua1 = 3.989089634e-09 lua1 = -7.227073177e-16   ub1 = -4.632061037e-18 lub1 = 9.614603776e-25 wub1 = -5.877471754e-39   uc1 = -1.636467021e-10 luc1 = 7.779412089e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.5 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.903453451e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.917847848e-8   k1 = 3.085216440e-01 lk1 = 5.473565751e-8   k2 = 4.751743479e-03 lk2 = -1.488387669e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.102284893e+05 lvsat = 8.563871006e-3   ua = -1.694891786e-09 lua = -4.934109040e-17   ub = 2.753384219e-18 lub = 1.966037765e-26   uc = 7.295344036e-11 luc = -3.761463173e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.510098374e-02 lu0 = -4.352250051e-11   a0 = 1.333329778e+00 la0 = 5.644842443e-8   keta = -1.316929513e-02 lketa = 1.720119165e-9   a1 = 0.0   a2 = 0.38689047   ags = 2.402114010e+00 lags = -4.844943852e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.181877789e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.707009101e-9   nfactor = {2.061400887e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.649358879e-08 wnfactor = -3.388131789e-21   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -4.638664827e-03 leta0 = 2.099778659e-09 weta0 = -1.990403349e-24 peta0 = 8.597351272e-31   etab = 2.191282287e-02 letab = -9.926128151e-09 wetab = 1.209751646e-23 petab = -2.761013168e-30   dsub = 1.588821784e+00 ldsub = -2.659678555e-7   voffl = 0.0   minv = 0.0   pclm = 6.274339786e-01 lpclm = -4.987795901e-08 wpclm = -8.470329473e-22   pdiblc1 = 0.39   pdiblc2 = 7.760005620e-03 lpdiblc2 = 1.246675661e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.021198007e-03 lalpha0 = 9.851108341e-10 walpha0 = 8.271806126e-25 palpha0 = 4.437342592e-31   alpha1 = 0.0   beta0 = 1.882254688e+01 lbeta0 = 2.510258883e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.549086746e-01 lkt1 = -3.618675627e-9   kt2 = -2.800928594e-02 lkt2 = 1.283846348e-9   at = 8.582104642e+04 lat = -6.172884838e-3   ute = -4.899828300e-01 lute = -2.374186476e-7   ua1 = 3.921070339e-09 lua1 = -6.919833421e-16   ub1 = -3.957051323e-18 lub1 = 6.565618647e-25   uc1 = 4.498102275e-11 luc1 = -1.644197929e-17 puc1 = -8.816207631e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.6 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.948835671e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.026331517e-8   k1 = 3.567334157e-01 lk1 = 4.501158422e-8   k2 = -2.989071599e-02 lk2 = -7.896665828e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.470853184e+05 lvsat = 1.130032860e-3   ua = -1.102729397e-09 lua = -1.687772834e-16   ub = 3.088596943e-18 lub = -4.795035268e-26   uc = 7.869818671e-11 luc = -4.920149789e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.577484904e-02 lu0 = -4.213337762e-9   a0 = 4.648205343e+00 la0 = -6.121454026e-7   keta = 2.073280580e-01 lketa = -4.275309447e-08 wketa = -5.293955920e-23 pketa = 1.735493991e-29   a1 = 0.0   a2 = 0.38689047   ags = -2.264777729e+00 lags = 4.567943440e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.555092897e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.234571230e-9   nfactor = {7.519402440e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.906052532e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.290661926e-01 leta0 = 2.719618888e-08 weta0 = -7.940933881e-23 peta0 = -9.466330863e-30   etab = -5.076770586e-02 letab = 4.733171092e-9   dsub = 1.728030840e-01 ldsub = 1.963603610e-8   voffl = 0.0   minv = 0.0   pclm = 8.162573993e-01 lpclm = -8.796269885e-8   pdiblc1 = -7.576278571e-01 lpdiblc1 = 2.314708006e-7   pdiblc2 = 1.437935621e-02 lpdiblc2 = -8.841425664e-11   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 7.038427000e-03 lalpha0 = -8.421702317e-10   alpha1 = 0.0   beta0 = 3.553786598e+01 lbeta0 = -8.611374045e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.962787643e-01 lkt1 = -1.544403539e-8   kt2 = -3.301492257e-02 lkt2 = 2.293458228e-09 wkt2 = -5.293955920e-23   at = 8.703207357e+03 lat = 9.381397712e-3   ute = -1.221594629e+00 lute = -8.985620589e-8   ua1 = 1.378170368e-09 lua1 = -1.790931325e-16 wua1 = 1.577721810e-30   ub1 = -1.794635110e-18 lub1 = 2.204133267e-25   uc1 = -1.088225635e-10 luc1 = 1.457943503e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.7 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.935173720e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = -1.057489410e-8   k1 = 9.509947867e-01 lk1 = -3.324966703e-8   k2 = -2.267425973e-01 lk2 = 1.802774268e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.648965162e+05 lvsat = -1.215612827e-3   ua = -3.245751423e-09 lua = 1.134480023e-16   ub = 3.834955308e-18 lub = -1.462420176e-25   uc = 1.584401315e-10 luc = -1.542176521e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.151152862e-02 lu0 = 2.989702203e-10   a0 = 0.0   keta = 1.041168850e-01 lketa = -2.916069905e-8   a1 = 0.0   a2 = 0.38689047   ags = 1.043460883e+00 lags = 2.111585997e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.128084382e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.611082588e-9   nfactor = {1.295907430e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.189674947e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 6.952563100e-02 leta0 = 1.042638666e-9   etab = -6.508939773e-02 letab = 6.619266302e-9   dsub = 5.317546079e-01 ldsub = -2.763608485e-8   voffl = 0.0   minv = 0.0   pclm = 9.866894167e-02 lpclm = 6.540113077e-9   pdiblc1 = 3.086130789e+00 lpdiblc1 = -2.747329943e-7   pdiblc2 = 5.490905128e-02 lpdiblc2 = -5.425972449e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.486389796e-03 lalpha0 = -1.109946920e-10   alpha1 = 0.0   beta0 = 3.080910576e+01 lbeta0 = -2.383833271e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.986686317e-01 lkt1 = -1.959801803e-9   kt2 = 1.413561800e-02 lkt2 = -3.916032213e-9   at = 6.702373500e+04 lat = 1.700875824e-3   ute = -2.660849783e+00 lute = 9.968650172e-8   ua1 = -1.957732867e-09 lua1 = 2.602286440e-16 wua1 = 5.916456789e-31 pua1 = 3.526483052e-38   ub1 = 1.950353760e-18 lub1 = -2.727829826e-25 wub1 = -7.346839693e-40 pub1 = 1.751623080e-46   uc1 = 4.573332750e-12 luc1 = -3.542375240e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.8 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.948091846e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.600903740e-7   k1 = 6.578690425e-01 wk1 = -1.298880553e-6   k2 = -9.751470123e-02 wk2 = 4.434986054e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -5.043492431e+04 wvsat = 1.479551909e+0   ua = -1.394124282e-09 wua = 6.473071250e-16   ub = 2.698968817e-18 wub = -8.264945878e-26   uc = 6.940459561e-11 wuc = 5.226628794e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.103021879e-02 wu0 = 7.567037210e-9   a0 = 2.047916618e+00 wa0 = -6.441541476e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.054006181e-01 wags = 3.435287679e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.070539010e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -5.975754807e-8   nfactor = {1.206922917e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.178851837e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 5.402215816e-01 wpclm = -2.379183129e-6   pdiblc1 = 0.39   pdiblc2 = 1.702582195e-04 wpdiblc2 = 3.235988547e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.150915353e-04 walpha0 = -9.143111569e-10   alpha1 = 0.0   beta0 = 1.855131594e+01 wbeta0 = -5.093268376e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.526313920e-01 wkt1 = -7.053236088e-9   kt2 = -3.373249145e-02 wkt2 = -4.828753937e-9   at = 1.018377413e+06 wat = -4.792312218e+0   ute = -7.694280164e-01 wute = -2.155758312e-6   ua1 = 2.053859631e-09 wua1 = 4.394708640e-15   ub1 = -2.972925169e-19 wub1 = -1.500711617e-23   uc1 = 8.327821538e-13 wuc1 = -1.402508868e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.9 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.948091846e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.600903740e-7   k1 = 6.578690425e-01 wk1 = -1.298880553e-6   k2 = -9.751470123e-02 wk2 = 4.434986054e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -5.043492431e+04 wvsat = 1.479551909e+0   ua = -1.394124282e-09 wua = 6.473071250e-16   ub = 2.698968817e-18 wub = -8.264945878e-26   uc = 6.940459561e-11 wuc = 5.226628794e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.103021879e-02 wu0 = 7.567037210e-9   a0 = 2.047916618e+00 wa0 = -6.441541476e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.054006181e-01 wags = 3.435287679e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.070539010e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -5.975754807e-8   nfactor = {1.206922917e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.178851837e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 5.402215816e-01 wpclm = -2.379183129e-6   pdiblc1 = 0.39   pdiblc2 = 1.702582195e-04 wpdiblc2 = 3.235988547e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.150915353e-04 walpha0 = -9.143111569e-10   alpha1 = 0.0   beta0 = 1.855131594e+01 wbeta0 = -5.093268376e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.526313920e-01 wkt1 = -7.053236088e-9   kt2 = -3.373249145e-02 wkt2 = -4.828753937e-9   at = 1.018377413e+06 wat = -4.792312218e+0   ute = -7.694280164e-01 wute = -2.155758312e-6   ua1 = 2.053859631e-09 wua1 = 4.394708640e-15   ub1 = -2.972925169e-19 wub1 = -1.500711617e-23   uc1 = 8.327821538e-13 wuc1 = -1.402508868e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.10 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.525924493e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.668276618e-07 wvth0 = 3.662074767e-07 pvth0 = -8.145119243e-13   k1 = 1.043642792e+00 lk1 = -1.524460197e-06 wk1 = -3.711772187e-06 pk1 = 9.535011802e-12   k2 = -2.324318590e-01 lk2 = 5.331514576e-07 wk2 = 1.285360044e-06 pk2 = -3.326779636e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.361573984e+05 lvsat = 3.387490723e-01 wvsat = 2.868217635e+00 pvsat = -5.487583409e-6   ua = -1.626157935e-09 lua = 9.169262272e-16 wua = 1.750072901e-15 pua = -4.357794004e-21   ub = 2.590227937e-18 lub = 4.297107919e-25 wub = 3.816804042e-25 pub = -1.834889998e-30   uc = 1.249389400e-10 luc = -2.194547912e-16 wuc = -4.021870879e-16 puc = 1.609974747e-21   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.498735124e-02 lu0 = 2.387956948e-08 wu0 = 3.531529099e-08 pu0 = -1.096526357e-13   a0 = 1.946138753e+00 la0 = 4.021950800e-07 wa0 = -2.116452637e-07 pa0 = -1.709143194e-12   keta = 1.006519294e-01 lketa = -3.977457260e-07 wketa = 5.553956970e-07 pketa = -2.194754399e-12   a1 = 0.0   a2 = 0.38689047   ags = -7.282625602e-01 lags = 4.875060613e-06 wags = 2.281702680e-06 pags = -7.659072156e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.695214666e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.943600195e-08 wvoff = -1.983006252e-07 pvoff = 5.474799854e-13   nfactor = {1.424787696e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.609351597e-07 wnfactor = -4.510381542e-06 pnfactor = 1.316518928e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.618558914e-06 lcit = 4.986469617e-11 wcit = 8.824208723e-11 pcit = -3.487058149e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378214013e-01 letab = 2.680094922e-7   dsub = 1.179574406e+00 ldsub = -2.448369081e-06 wdsub = -2.442240951e-06 pdsub = 9.650991356e-12   voffl = 0.0   minv = 0.0   pclm = 3.865810037e-01 lpclm = 6.071407036e-07 wpclm = -1.510175054e-06 ppclm = -3.434054865e-12   pdiblc1 = 0.39   pdiblc2 = -7.913245156e-03 lpdiblc2 = 3.194353987e-08 wpdiblc2 = 6.231630924e-08 ppdiblc2 = -1.183786500e-13   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.106215500e-04 lalpha0 = -3.775054814e-10 walpha0 = -1.865107628e-09 palpha0 = 3.757257662e-15   alpha1 = 0.0   beta0 = 1.592482568e+01 lbeta0 = 1.037908843e-05 wbeta0 = -1.043060867e-05 pbeta0 = 2.109154095e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.793420211e-01 lkt1 = 1.055522596e-07 wkt1 = 1.796670205e-07 pkt1 = -7.378615043e-13   kt2 = -1.800888339e-02 lkt2 = -6.213490333e-08 wkt2 = -1.473220764e-07 pkt2 = 5.630901499e-13   at = 1.979313845e+06 lat = -3.797327695e+00 wat = -9.589805071e+00 pat = 1.895822852e-5   ute = -5.413338221e-01 lute = -9.013586872e-07 wute = -3.126421272e-06 pute = 3.835763964e-12   ua1 = -6.864508227e-10 lua1 = 1.082887112e-14 wua1 = 1.966941394e-14 pua1 = -6.036097656e-20   ub1 = 5.337801999e-18 lub1 = -2.226817482e-23 wub1 = -4.538180743e-23 pub1 = 1.200315156e-28   uc1 = 2.356404479e-11 luc1 = -8.982701689e-17 wuc1 = -1.932667328e-16 puc1 = 2.095024536e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.11 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.365885512e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.892889600e-09 wvth0 = -6.595840021e-08 pvth0 = 2.894405689e-14   k1 = 1.107984551e-01 lk1 = 2.961674307e-07 wk1 = 2.225532567e-06 pk1 = -2.052796199e-12   k2 = 9.846654331e-02 lk2 = -1.126612996e-07 wk2 = -7.936687868e-07 pk2 = 7.308505373e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.869953906e+03 lvsat = 5.765160891e-02 wvsat = 8.369345356e-02 pvsat = -5.304148580e-8   ua = -8.827073103e-10 lua = -5.340626402e-16 wua = -5.173925089e-16 pua = 6.760689951e-23   ub = 2.698509633e-18 lub = 2.183779469e-25 wub = -3.725861836e-25 pub = -3.627916698e-31   uc = -8.353095905e-11 luc = 1.874148685e-16 wuc = 1.003684774e-15 puc = -1.133858336e-21   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.243251155e-02 lu0 = -1.016806267e-08 wu0 = -2.912354438e-08 pu0 = 1.611231708e-14   a0 = 2.488260506e+00 la0 = -6.558612341e-07 wa0 = -2.115549302e-06 pa0 = 2.006696798e-12   keta = 1.507962877e-01 lketa = -4.956122195e-07 wketa = -2.074813903e-06 pketa = 2.938612526e-12   a1 = 0.0   a2 = 0.38689047   ags = 9.730782217e-01 lags = 1.554562316e-06 wags = -5.897879400e-07 pags = -2.054798271e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.420930652e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.818225300e-08 wvoff = 1.752035249e-07 pvoff = -1.814861969e-13   nfactor = {-2.988476735e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.978141815e-06 wnfactor = 6.284644705e-06 pnfactor = -7.903409473e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 3.999559283e-05 lcit = -3.330513072e-11 wcit = -1.764841745e-10 pcit = 1.679591064e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 7.515109248e-04 leta0 = -4.908726144e-10 weta0 = -1.136827115e-09 peta0 = 2.218739796e-15   etab = -5.871773009e-04 letab = 1.701435022e-10 wetab = 3.259879720e-10 petab = -6.362290951e-16   dsub = 1.795012591e-01 ldsub = -4.965313211e-07 wdsub = -1.557476567e-06 pdsub = 7.924201131e-12   voffl = 0.0   minv = 0.0   pclm = 1.246153854e+00 lpclm = -1.070483330e-06 wpclm = -7.111228407e-06 ppclm = 7.497492959e-12   pdiblc1 = 0.39   pdiblc2 = 1.057540683e-02 lpdiblc2 = -4.140669762e-09 wpdiblc2 = -2.460461257e-08 ppdiblc2 = 5.126447846e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.593214078e-04 lalpha0 = -8.221375036e-11 walpha0 = 1.801528646e-10 palpha0 = -2.344670159e-16   alpha1 = 0.0   beta0 = 2.069229504e+01 lbeta0 = 1.074442309e-06 wbeta0 = 3.546397014e-06 pbeta0 = -6.187311154e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.145095509e-01 lkt1 = -2.098094835e-08 wkt1 = -2.534720368e-07 pkt1 = 1.074938281e-13   kt2 = -1.407521292e-01 lkt2 = 1.774224758e-07 wkt2 = 6.657841060e-07 pkt2 = -1.023845121e-12   at = 5.925004143e+02 lat = 6.453285934e-02 wat = 2.161569727e-01 pat = -1.800185702e-7   ute = -1.396674033e+00 lute = 7.680045259e-07 wute = 5.325516610e-07 pute = -3.305435214e-12   ua1 = 3.823005348e-09 lua1 = 2.027788056e-15 wua1 = -3.843286534e-15 pua1 = -1.447135661e-20   ub1 = -4.804233559e-18 lub1 = -2.474014733e-24 wub1 = 6.289804403e-24 pub1 = 1.918428913e-29   uc1 = 1.665354911e-10 luc1 = -3.688636738e-16 wuc1 = -1.093748950e-15 puc1 = 1.966969095e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.12 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.488489554e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.775275756e-09 wvth0 = -4.444667206e-08 pvth0 = 8.471452763e-15   k1 = 4.484269207e-01 lk1 = -2.515189183e-08 wk1 = -1.030060928e-07 pk1 = 1.632624011e-13   k2 = -2.709125547e-02 lk2 = 6.831429702e-09 wk2 = 5.358554291e-08 pk2 = -7.547717207e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.344155490e+05 lvsat = -6.278120125e-02 wvsat = -7.918192205e-01 pvsat = 7.801795485e-7   ua = -6.830447064e-10 lua = -7.240805419e-16 wua = -3.894260229e-15 pua = 3.281355025e-21   ub = 2.572845460e-18 lub = 3.379719121e-25 wub = 1.876627217e-24 pub = -2.503356817e-30   uc = 1.369101149e-10 luc = -2.237779939e-17 wuc = -2.136400696e-16 puc = 2.466363112e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.992521534e-02 lu0 = -7.781881411e-09 wu0 = -3.778690638e-08 pu0 = 2.435719537e-14   a0 = 2.356513468e+00 la0 = -5.304782371e-07 wa0 = -1.758220997e-06 pa0 = 1.666629237e-12   keta = -6.738728369e-01 lketa = 2.892212631e-07 wketa = 1.775102443e-06 pketa = -7.253336113e-13   a1 = 0.0   a2 = 0.38689047   ags = 7.755633402e-01 lags = 1.742536241e-06 wags = 1.563959532e-05 pags = -1.750022117e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.109258873e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.479394317e-09 wvoff = -2.818046813e-08 pvoff = 1.207333231e-14   nfactor = {2.570064511e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.962169142e-07 wnfactor = -7.941906823e-06 pnfactor = 5.635928484e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.162760515e-04 leta0 = -1.718312220e-10 weta0 = 2.437034305e-09 peta0 = -1.182486248e-15   etab = -7.223706044e-04 letab = 2.988062932e-10 wetab = -6.417559158e-10 petab = 2.847679243e-16   dsub = -1.554791741e+00 ldsub = 1.153986655e-06 wdsub = 1.288391694e-05 pdsub = -5.819600862e-12   voffl = 0.0   minv = 0.0   pclm = -5.453006658e-01 lpclm = 6.344349789e-07 wpclm = 3.621716801e-06 ppclm = -2.716997331e-12   pdiblc1 = 0.39   pdiblc2 = 8.689662698e-04 lpdiblc2 = 5.096901185e-09 wpdiblc2 = 6.601260137e-08 ppdiblc2 = -3.497547096e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -9.911261092e-05 lalpha0 = 1.637366131e-10 walpha0 = 5.288253512e-10 palpha0 = -5.662968780e-16   alpha1 = 0.0   beta0 = 1.848143833e+01 lbeta0 = 3.178503594e-06 wbeta0 = 1.566744672e-06 pbeta0 = -4.303285918e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.189058275e-01 lkt1 = -1.679703388e-08 wkt1 = -2.243361439e-07 pkt1 = 7.976534456e-14   kt2 = 8.804468444e-02 lkt2 = -4.032230776e-08 wkt2 = -6.291861581e-07 pkt2 = 2.085716047e-13   at = 1.386723905e+04 lat = 5.189935695e-02 wat = 4.090328654e-01 pat = -3.635775929e-7   ute = -2.726768496e-01 lute = -3.016979736e-07 wute = -5.123414703e-06 pute = 2.077319694e-12   ua1 = 9.209702971e-09 lua1 = -3.098705138e-15 wua1 = -3.650795789e-14 pua1 = 1.661544780e-20   ub1 = -1.194894071e-17 lub1 = 4.325567342e-24 wub1 = 5.116723225e-23 pub1 = -2.352533456e-29   uc1 = -5.094186612e-10 luc1 = 2.744385132e-16 wuc1 = 2.417997141e-15 puc1 = -1.375142101e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.13 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.892424914e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.702083400e-08 wvth0 = 7.712300090e-09 pvth0 = -1.508849416e-14   k1 = 2.862539876e-01 lk1 = 4.810081120e-08 wk1 = 1.557186119e-07 pk1 = 4.639774565e-14   k2 = 2.068321615e-02 lk2 = -1.474806026e-08 wk2 = -1.114094256e-07 pk2 = -9.497697622e-16   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.345286527e+05 lvsat = 5.869954997e-02 wvsat = 1.711596485e+00 pvsat = -3.506008084e-7   ua = -2.053631787e-09 lua = -1.049932105e-16 wua = 2.508683178e-15 pua = 3.891775022e-22   ub = 3.302274752e-18 lub = 8.492347990e-27 wub = -3.838413453e-24 pub = 7.809847812e-32   uc = 1.301661585e-10 luc = -1.933158801e-17 wuc = -4.000908266e-16 puc = 1.088825058e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.589952555e-02 lu0 = -1.446547459e-09 wu0 = -5.584234844e-09 pu0 = 9.811409652e-15   a0 = 4.860584913e-01 la0 = 3.143969238e-07 wa0 = 5.925001999e-06 pa0 = -1.803844174e-12   keta = -1.210546937e-01 lketa = 3.951607185e-08 wketa = 7.544469075e-07 pketa = -2.643086090e-13   a1 = 0.0   a2 = 0.38689047   ags = 8.371417296e+00 lags = -1.688473011e-06 wags = -4.174357665e-05 pags = 8.419470692e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.222475104e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.634526199e-09 wvoff = 2.838986468e-08 pvoff = -1.347920417e-14   nfactor = {1.276744839e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.796911543e-08 wnfactor = 5.487131135e-06 pnfactor = -4.299008168e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -9.154619865e-03 leta0 = 4.151295004e-09 weta0 = 3.158026062e-08 peta0 = -1.434633586e-14   etab = -3.847765836e-02 letab = 1.735268100e-08 wetab = 4.223130508e-07 petab = -1.907618035e-13   dsub = 1.733502234e+00 ldsub = -3.313192916e-07 wdsub = -1.011756178e-06 pdsub = 4.570052067e-13   voffl = 0.0   minv = 0.0   pclm = 1.271559315e+00 lpclm = -1.862315903e-07 wpclm = -4.504394245e-06 ppclm = 9.535263979e-13   pdiblc1 = 0.39   pdiblc2 = 1.274462754e-02 lpdiblc2 = -2.672756333e-10 wpdiblc2 = -3.485766048e-08 ppdiblc2 = 1.058712196e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.960376926e-03 lalpha0 = 1.907850398e-09 walpha0 = 1.356075575e-08 palpha0 = -6.452754679e-15   alpha1 = 0.0   beta0 = 1.926987033e+01 lbeta0 = 2.822372798e-06 wbeta0 = -3.128150844e-06 pbeta0 = -2.182625088e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.858416623e-01 lkt1 = -3.173195197e-08 wkt1 = -4.829883793e-07 pkt1 = 1.965972660e-13   kt2 = 6.284512546e-03 lkt2 = -3.391646913e-09 wkt2 = -2.398179046e-07 pkt2 = 3.269591139e-14   at = 1.744222187e+05 lat = -2.062252456e-02 wat = -6.195915415e-01 pat = 1.010469086e-7   ute = 1.372414829e+00 lute = -1.044777659e-06 wute = -1.302382132e-05 pute = 5.645893862e-12   ua1 = 8.120110698e-09 lua1 = -2.606541756e-15 wua1 = -2.936405720e-14 pua1 = 1.338858357e-20   ub1 = -7.195366116e-18 lub1 = 2.178401464e-24 wub1 = 2.264566488e-23 pub1 = -1.064228519e-29   uc1 = 2.830603095e-10 luc1 = -8.352027551e-17 wuc1 = -1.664897976e-15 puc1 = 4.690812085e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.14 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.821698758e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.576382279e-08 wvth0 = 8.890735207e-08 pvth0 = -3.146513017e-14   k1 = 2.226029659e-01 lk1 = 6.093890402e-08 wk1 = 9.379796005e-07 pk1 = -1.113803844e-13   k2 = 2.822936529e-02 lk2 = -1.627008081e-08 wk2 = -4.064360532e-07 pk2 = 5.855562589e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.666739337e+05 lvsat = -2.051505698e-03 wvsat = -1.369839700e-01 pvsat = 2.224862639e-8   ua = -3.014333955e-09 lua = 8.877561314e-17 wua = 1.336792713e-14 pua = -1.801077708e-21   ub = 4.771855341e-18 lub = -2.879147090e-25 wub = -1.177109331e-23 pub = 1.678080342e-30   uc = -6.162851219e-12 luc = 8.165291605e-18 wuc = 5.934366327e-16 puc = -9.150701509e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.024827622e-02 lu0 = -2.323668726e-09 wu0 = 1.085779447e-07 pu0 = -1.321453116e-14   a0 = 5.891892731e+00 la0 = -7.759328132e-07 wa0 = -8.697155655e-06 pa0 = 1.145371914e-12   keta = 5.965207483e-01 lketa = -1.052153069e-07 wketa = -2.721640051e-06 pketa = 4.368007501e-13   a1 = 0.0   a2 = 0.38689047   ags = -2.322677388e+00 lags = 4.684724158e-07 wags = 4.048946347e-07 pags = -8.166522334e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.636574168e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.198669727e-08 wvoff = 5.698017844e-08 pvoff = -1.924572750e-14   nfactor = {-3.720992927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.205327325e-07 wnfactor = 7.860453442e-06 pnfactor = -9.085880596e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.486488789e-07 lcit = 8.978152644e-13 wcit = 3.112847644e-11 pcit = -6.278458056e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -4.696315241e-02 leta0 = 1.177708679e-08 weta0 = -5.741498443e-07 peta0 = 1.078263976e-13   etab = 1.543946902e-01 letab = -2.154870735e-08 wetab = -1.434708842e-06 petab = 1.837902272e-13   dsub = -3.629953708e-01 ldsub = 9.153379279e-08 wdsub = 3.746860026e-06 pdsub = -5.027838885e-13   voffl = 0.0   minv = 0.0   pclm = 6.702476199e-01 lpclm = -6.495002791e-08 wpclm = 1.021052228e-06 ppclm = -1.609285284e-13   pdiblc1 = -7.576349608e-01 lpdiblc1 = 2.314722334e-07 wpdiblc1 = 4.967614846e-11 ppdiblc1 = -1.001943076e-17   pdiblc2 = -1.026080681e-02 lpdiblc2 = 4.372805448e-09 wpdiblc2 = 1.723096456e-07 ppdiblc2 = -3.119748784e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.867914251e-02 lalpha0 = -2.658427474e-09 walpha0 = -8.140398915e-08 palpha0 = 1.270115954e-14   alpha1 = 0.0   beta0 = 4.805262809e+01 lbeta0 = -2.982965527e-06 wbeta0 = -8.751623197e-05 pbeta0 = 1.483802893e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.765575429e-01 lkt1 = 6.734487561e-09 wkt1 = 1.260696710e-06 pkt1 = -1.550952981e-13   kt2 = -7.690194233e-02 lkt2 = 1.338664510e-08 wkt2 = 3.069036847e-07 pkt2 = -7.757509955e-14   at = 7.265450781e+04 lat = -9.648612119e-05 wat = -4.472140021e-01 pat = 6.627922076e-8   ute = -5.856423953e+00 lute = 4.132429788e-07 wute = 3.241154686e-05 pute = -3.518192723e-12   ua1 = -1.256073034e-08 lua1 = 1.564680477e-15 wua1 = 9.747529020e-14 pua1 = -1.219427860e-20   ub1 = 1.037877363e-17 lub1 = -1.366214653e-24 wub1 = -8.512913427e-23 pub1 = 1.109535292e-29   uc1 = -3.902566868e-10 luc1 = 5.228439607e-17 wuc1 = 1.968080082e-15 puc1 = -2.636723007e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.15 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.210993591e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.455164109e-08 wvth0 = -8.921859390e-07 pvth0 = 9.773995079e-14   k1 = 1.419447798e+00 lk1 = -9.667957615e-08 wk1 = -3.275910647e-06 pk1 = 4.435678917e-13   k2 = -3.748380569e-01 lk2 = 3.681188336e-08 wk2 = 1.035637473e-06 pk2 = -1.313582471e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.065497604e+04 lvsat = 9.276760928e-03 wvsat = 5.891044598e-01 pvsat = -7.337358936e-8   ua = -6.145064839e-09 lua = 5.010772169e-16 wua = 2.027501469e-14 pua = -2.710706603e-21   ub = 7.741532788e-18 lub = -6.790063803e-25 wub = -2.731885258e-23 pub = 3.725642499e-30   uc = 3.434627704e-10 luc = -3.787865464e-17 wuc = -1.293870715e-15 puc = 1.570419261e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 5.089632512e-03 lu0 = 9.895988577e-10 wu0 = 4.490857634e-08 pu0 = -4.829593686e-15   a0 = 0.0   keta = 4.455050342e-01 lketa = -8.532729246e-08 wketa = -2.387340983e-06 pketa = 3.927752344e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.184696779e+00 lags = 6.568774878e-09 wags = -9.876682665e-07 pags = 1.017283479e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-3.545064694e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.712056326e-08 wvoff = 1.690204000e-06 pvoff = -2.343331387e-13   nfactor = {-1.722945935e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.984324811e-07 wnfactor = 2.111096234e-05 pnfactor = -2.653613828e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.538648595e-05 lcit = -1.056253689e-12 wcit = -7.263311170e-11 pcit = 7.386424295e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.458389392e-01 leta0 = 3.796803353e-08 weta0 = 2.205357054e-06 peta0 = -2.582207633e-13   etab = -1.443454137e-01 letab = 1.779387064e-08 wetab = 5.542404902e-07 petab = -7.814445511e-14   dsub = 5.762805813e-01 ldsub = -3.216415372e-08 wdsub = -3.113719132e-07 pdsub = 3.166496671e-14   voffl = 0.0   minv = 0.0   pclm = 1.149510897e+00 lpclm = -1.280666052e-07 wpclm = -7.348579830e-06 ppclm = 9.413101655e-13   pdiblc1 = 7.493555756e+00 lpdiblc1 = -8.551683280e-07 wpdiblc1 = -3.082129909e-05 ppdiblc1 = 4.059007506e-12   pdiblc2 = 1.075157751e-01 lpdiblc2 = -1.113778150e-08 wpdiblc2 = -3.678809237e-07 ppdiblc2 = 3.994290918e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.748625037e-03 lalpha0 = 5.585873727e-10 walpha0 = 5.059474812e-08 palpha0 = -4.682414162e-15   alpha1 = 0.0   beta0 = 2.119235472e+01 lbeta0 = 5.543981745e-07 wbeta0 = 6.725032474e-05 pbeta0 = -5.543952752e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 1.417939780e-02 lkt1 = -4.472361385e-08 wkt1 = -2.187758784e-06 pkt1 = 2.990490482e-13   kt2 = 3.001868264e-01 lkt2 = -3.627406030e-08 wkt2 = -2.000367543e-06 pkt2 = 2.262809847e-13   at = -4.945501850e+04 lat = 1.598472795e-02 wat = 8.145405824e-01 pat = -9.988754925e-8   ute = -3.988346659e+00 lute = 1.672265396e-07 wute = 9.283238753e-06 pute = -4.723101868e-13   ua1 = -5.713001815e-09 lua1 = 6.628688687e-16 wua1 = 2.626074597e-14 pua1 = -2.815679197e-21   ub1 = 4.847345191e-18 lub1 = -6.377531841e-25 wub1 = -2.025877696e-23 pub1 = 2.552251218e-30   uc1 = -2.099203598e-10 luc1 = 2.853500348e-17 wuc1 = 1.499962972e-15 puc1 = -2.020236179e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.16 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.426554+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40031   k2 = -0.009571991   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 242950.0   ua = -1.26576775e-9   ub = 2.68258e-18   uc = 7.0441e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03253071   a0 = 1.9201853   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.57352   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.97316474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.068446   pdiblc1 = 0.39   pdiblc2 = 0.006587   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.3789948e-5   alpha1 = 0.0   beta0 = 17.541356   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25403   kt2 = -0.03469   at = 68095.0   ute = -1.1969   ua1 = 2.9253e-9   ub1 = -3.2731e-18   uc1 = -2.6978e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.17 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.426554+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40031   k2 = -0.009571991   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 242950.0   ua = -1.26576775e-9   ub = 2.68258e-18   uc = 7.0441e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03253071   a0 = 1.9201853   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.57352   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.97316474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.068446   pdiblc1 = 0.39   pdiblc2 = 0.006587   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.3789948e-5   alpha1 = 0.0   beta0 = 17.541356   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25403   kt2 = -0.03469   at = 68095.0   ute = -1.1969   ua1 = 2.9253e-9   ub1 = -3.2731e-18   uc1 = -2.6978e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.18 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.252088625e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.315573012e-9   k1 = 3.076240044e-01 lk1 = 3.662667852e-7   k2 = 2.244615977e-02 lk2 = -1.265259663e-07 pk2 = 3.231174268e-27   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.325903481e+05 lvsat = -7.494008152e-1   ua = -1.279130567e-09 lua = 5.280577528e-17   ub = 2.665912525e-18 lub = 6.586477881e-26   uc = 4.518801839e-11 luc = 9.979208114e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.199012952e-02 lu0 = 2.136209184e-9   a0 = 1.904170959e+00 la0 = 6.328378955e-8   keta = 2.107830600e-01 lketa = -8.329503643e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.758166784e-01 lags = 3.356319505e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.262737910e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.912549774e-8   nfactor = {5.304101896e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.749630943e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.487923750e-05 lcit = -1.928125843e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378214013e-01 letab = 2.680094922e-7   dsub = 6.952948933e-01 ldsub = -5.346441536e-7   voffl = 0.0   minv = 0.0   pclm = 8.712372115e-02 lpclm = -7.380865728e-8   pdiblc1 = 0.39   pdiblc2 = 4.443648551e-03 lpdiblc2 = 8.469871204e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.921641048e-05 lalpha0 = 3.675327618e-10   alpha1 = 0.0   beta0 = 1.385650802e+01 lbeta0 = 1.456139532e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.437152919e-01 lkt1 = -4.076058033e-8   kt2 = -4.722183359e-02 lkt2 = 4.952198416e-8   at = 7.772173559e+04 lat = -3.804192289e-2   ute = -1.161281566e+00 lute = -1.407531866e-7   ua1 = 3.213858106e-09 lua1 = -1.140293624e-15   ub1 = -3.661096966e-18 lub1 = 1.533245671e-24   uc1 = -1.475941345e-11 luc1 = -4.828412737e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.19 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.235094560e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.632296166e-9   k1 = 5.521061915e-01 lk1 = -1.108878769e-7   k2 = -5.891249529e-02 lk2 = 3.226131398e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.446578768e+04 lvsat = 4.713384863e-2   ua = -9.853026712e-10 lua = -5.206566590e-16   ub = 2.624628366e-18 lub = 1.464388645e-25   uc = 1.154927992e-10 luc = -3.742140796e-17 wuc = -1.262177448e-29   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.665751385e-02 lu0 = -6.973101482e-9   a0 = 2.068761691e+00 la0 = -2.579471191e-07 wa0 = -2.168404345e-19   keta = -2.606249786e-01 lketa = 8.709434751e-8   a1 = 0.0   a2 = 0.38689047   ags = 8.561273468e-01 lags = 1.147110011e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.073514163e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.805206339e-9   nfactor = {1.216316870e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.109503045e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.260859600e-04 leta0 = -5.091183760e-11   etab = -5.225361376e-04 letab = 4.398366707e-11   dsub = -1.293355867e-01 ldsub = 1.074783031e-6   voffl = 0.0   minv = 0.0   pclm = -1.639536224e-01 lpclm = 4.162177387e-07 wpclm = -6.776263578e-21 ppclm = 6.462348536e-27   pdiblc1 = 0.39   pdiblc2 = 5.696482098e-03 lpdiblc2 = 6.024722235e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.950444766e-04 lalpha0 = -1.287069402e-10   alpha1 = 0.0   beta0 = 2.139552108e+01 lbeta0 = -1.524587575e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.647713051e-01 lkt1 = 3.343353071e-10   kt2 = -8.731739510e-03 lkt2 = -2.559894002e-8   at = 4.345493513e+04 lat = 2.883642024e-2   ute = -1.291072717e+00 lute = 1.125595534e-7   ua1 = 3.060908174e-09 lua1 = -8.417820067e-16   ub1 = -3.557008789e-18 lub1 = 1.330097297e-24   uc1 = -5.034737131e-11 luc1 = 2.117271203e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.20 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.400354873e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.095445185e-9   k1 = 4.280015240e-01 lk1 = 7.221914667e-9   k2 = -1.646561243e-02 lk2 = -8.135172203e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.259673333e+04 lvsat = 9.192301456e-2   ua = -1.455249612e-09 lua = -7.341050466e-17   ub = 2.944967675e-18 lub = -1.584264542e-25   uc = 9.454676469e-11 luc = -1.748717169e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.243233280e-02 lu0 = -2.952017803e-9   a0 = 2.007870389e+00 la0 = -1.999971707e-7   keta = -3.218822829e-01 lketa = 1.453926178e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.876787069e+00 lags = -1.727636744e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.165138795e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.146640901e-10   nfactor = {9.952392426e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.213487771e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.995231701e-04 leta0 = -4.063100777e-10   etab = -8.496263699e-04 letab = 3.552738057e-10   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 1.728607608e-01 lpclm = 9.567317430e-8   pdiblc1 = 0.39   pdiblc2 = 1.395880918e-02 lpdiblc2 = -1.838493134e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 5.749803653e-06 lalpha0 = 5.144385357e-11   alpha1 = 0.0   beta0 = 1.879211297e+01 lbeta0 = 2.325191719e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.633901354e-01 lkt1 = -9.801169905e-10   kt2 = -3.671858495e-02 lkt2 = 1.036000854e-9   at = 9.497563110e+04 lat = -2.019556851e-2   ute = -1.288614598e+00 lute = 1.102201738e-7   ua1 = 1.970427080e-09 lua1 = 1.960233981e-16   ub1 = -1.802831967e-18 lub1 = -3.393440142e-25   uc1 = -2.994652916e-11 luc1 = 1.757332569e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.21 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.053454965e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.440823502e-07 wvth0 = 1.943720201e-06 pvth0 = -8.779686963e-13   k1 = 3.171319128e-01 lk1 = 5.730116370e-8   k2 = 3.210682617e-02 lk2 = -3.007509986e-08 wk2 = -1.690191479e-07 pk2 = 7.634510403e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.111712036e+05 lvsat = 3.150070631e-02 wvsat = 4.725222814e-01 pvsat = -2.134359519e-7   ua = -4.659794248e-09 lua = 1.374066285e-15 wua = 1.565166472e-14 pua = -7.069778694e-21   ub = 5.854005305e-18 lub = -1.472424206e-24 wub = -1.670689270e-23 pub = 7.546419898e-30   uc = 5.083091101e-11 luc = 2.259060844e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 6.869540392e-04 lu0 = 1.138721106e-08 wu0 = 1.215637718e-07 pu0 = -5.490974790e-14   a0 = 1.660945464e+00 la0 = -4.329291686e-8   keta = 2.854691715e-02 lketa = -1.289449974e-8   a1 = 0.0   a2 = 0.38689047   ags = 9.395436678e-02 lags = -1.895012601e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.166179963e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.616931123e-10   nfactor = {-8.537344970e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.927169403e-06 wnfactor = 5.497997860e-05 pnfactor = -2.483418143e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.892472934e-03 leta0 = 1.306515692e-9   etab = 4.526410273e-02 letab = -2.047406706e-08 wetab = 1.389663429e-21 petab = 7.415292509e-28   dsub = 1.532877972e+00 ldsub = -2.406983156e-7   voffl = 0.0   minv = 0.0   pclm = 3.783690482e-01 lpclm = 2.846108423e-9   pdiblc1 = 0.39   pdiblc2 = 5.832594228e-03 lpdiblc2 = 1.832077527e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.271372724e-03 lalpha0 = 6.283137138e-10 walpha0 = 5.293955920e-23 palpha0 = -1.893266173e-29   alpha1 = 0.0   beta0 = 1.864957963e+01 lbeta0 = 2.389573318e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.816149220e-01 lkt1 = 7.251927993e-9   kt2 = -4.126972152e-02 lkt2 = 3.091726487e-9   at = 5.156149546e+04 lat = -5.856205168e-4   ute = -1.210118985e+00 lute = 7.476409784e-8   ua1 = 2.297420972e-09 lua1 = 4.832189205e-17   ub1 = -2.704887182e-18 lub1 = 6.810981617e-26   uc1 = -4.707745968e-11 luc1 = 9.495288230e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.22 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.976322057e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.332842671e-07 wvth0 = -6.941857862e-06 pvth0 = 9.142079711e-13   k1 = 4.085978421e-01 lk1 = 3.885294308e-8   k2 = -1.720617026e-01 lk2 = 1.110467156e-08 wk2 = 6.036398140e-07 pk2 = -7.949634531e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.741463325e+05 lvsat = -4.170956233e-02 wvsat = -1.687579576e+00 pvsat = 2.222457923e-7   ua = 1.072078012e-08 lua = -1.728118663e-15 wua = -5.589880256e-14 pua = 7.361592803e-21   ub = -9.393919120e-18 lub = 1.603005911e-24 wub = 5.966747393e-23 pub = -7.857907979e-30   uc = 1.115115342e-10 luc = -9.979917453e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.378687338e-01 lu0 = -1.628166802e-08 wu0 = -4.341563278e-07 pu0 = 5.717621759e-14   a0 = 4.167306836e+00 la0 = -5.488134737e-7   keta = 5.683832440e-02 lketa = -1.860073513e-8   a1 = 0.0   a2 = 0.38689047   ags = -2.242389579e+00 lags = 4.522787660e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.523586409e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.170402438e-9   nfactor = {4.012282438e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.887343454e-06 wnfactor = -1.963570664e-04 pnfactor = 2.585924386e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 6.721210755e-06 lcit = -3.471596032e-13   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.608131009e-01 leta0 = 3.315831669e-08 weta0 = -5.929230631e-21   etab = -1.300981638e-01 letab = 1.489562528e-8   dsub = 3.799810930e-01 ldsub = -8.164779595e-9   voffl = 0.0   minv = 0.0   pclm = 8.727152243e-01 lpclm = -9.686104356e-8   pdiblc1 = -7.576251104e-01 lpdiblc1 = 2.314702466e-07 ppdiblc1 = -1.292469707e-26   pdiblc2 = 2.390700579e-02 lpdiblc2 = -1.813440912e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.537293709e-03 lalpha0 = -1.398752624e-10   alpha1 = 0.0   beta0 = 3.069876376e+01 lbeta0 = -4.068687485e-8   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.265700929e-01 lkt1 = -2.401983882e-8   kt2 = -1.604506143e-02 lkt2 = -1.995961330e-9   at = -1.602493993e+04 lat = 1.304622557e-2   ute = 5.705619243e-01 lute = -2.843903381e-7   ua1 = 6.767946451e-09 lua1 = -8.533607445e-16   ub1 = -6.501745711e-18 lub1 = 8.339171973e-25   uc1 = 0.0   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.23 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-6.078483166e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.070380502e-07 wvth0 = 4.296838348e-06 pvth0 = -5.658721262e-13   k1 = 7.698573433e-01 lk1 = -8.723126930e-9   k2 = -2.551217007e-01 lk2 = 2.204325800e-08 wk2 = 4.319030997e-07 pk2 = -5.687947871e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.143958949e+05 lvsat = -7.501728447e-03 wvsat = -8.535634381e-02 pvsat = 1.124100370e-8   ua = 7.445422114e-09 lua = -1.296770390e-15 wua = -4.826235463e-14 pua = 6.355910793e-21   ub = -1.762408783e-17 lub = 2.686877979e-24 wub = 1.006009868e-22 pub = -1.324864696e-29   uc = 8.689714433e-11 luc = -6.738325378e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 6.958504638e-02 lu0 = -7.289047799e-09 wu0 = -2.803443756e-07 pu0 = 3.691995255e-14   a0 = 0.0   keta = -2.788819345e-02 lketa = -7.442676360e-9   a1 = 0.0   a2 = 0.38689047   ags = 9.888489833e-01 lags = 2.674080364e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.935069032e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.346079620e-9   nfactor = {-3.067706069e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.436647410e-06 wnfactor = 1.671277212e-04 pnfactor = -2.200988524e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.838415715e-07 lcit = 4.084232314e-13   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.914681323e-01 leta0 = -1.323536032e-8   etab = -3.444335265e-02 letab = 2.298364930e-9   dsub = 5.145376816e-01 ldsub = -2.588520953e-8   voffl = 0.0   minv = 0.0   pclm = -3.076617267e-01 lpclm = 5.858869899e-8   pdiblc1 = 1.381905028e+00 lpdiblc1 = -5.029517490e-8   pdiblc2 = 3.456752883e-02 lpdiblc2 = -3.217378495e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.283964061e-03 lalpha0 = -3.699030145e-10   alpha1 = 0.0   beta0 = 3.452762962e+01 lbeta0 = -5.449293644e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.196380583e-01 lkt1 = 1.457574689e-8   kt2 = -9.647224083e-02 lkt2 = 8.595896062e-9   at = 1.120627530e+05 lat = -3.822283151e-3   ute = -2.147544533e+00 lute = 7.357069182e-8   ua1 = -5.056772717e-10 lua1 = 1.045391317e-16   ub1 = 8.301696467e-19 lub1 = -1.316593958e-25   uc1 = 8.751193733e-11 luc1 = -1.152488459e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.24 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.201373184e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.203874782e-8   k1 = 2.437293817e-01 wk1 = 7.818132904e-7   k2 = 5.099082976e-02 wk2 = -3.023925866e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.533532193e+05 wvsat = -5.512476901e-1   ua = -1.513984172e-09 wua = 1.239354524e-15   ub = 2.952053795e-18 wub = -1.345493439e-24   uc = 7.260003938e-11 wuc = -1.078016999e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.171789723e-02 wu0 = 4.058406654e-9   a0 = 2.279338622e+00 wa0 = -1.793266905e-6   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 6.229599982e-01 wags = -2.468558888e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.250892197e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 3.088599517e-8   nfactor = {5.552014819e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.086907266e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.754532663e-05 wcit = -3.767411769e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.300775800e-01 wpclm = 9.912361758e-7   pdiblc1 = 0.39   pdiblc2 = 6.399121367e-03 wpdiblc2 = 9.380855305e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.619336596e-05 walpha0 = 3.793003797e-11   alpha1 = 0.0   beta0 = 1.715745884e+01 wbeta0 = 1.916813899e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.513589544e-01 wkt1 = -1.333663766e-8   kt2 = -3.455418412e-02 wkt2 = -6.781341185e-10   at = -3.097523218e+05 wat = 1.886606792e+0   ute = -1.100168913e+00 wute = -4.829821888e-7   ua1 = 4.193518501e-09 wua1 = -6.332265702e-15   ub1 = -5.060436973e-18 wub1 = 8.924244999e-24   uc1 = 2.967892342e-12 wuc1 = -1.495210383e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.25 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.201373184e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.203874782e-8   k1 = 2.437293817e-01 wk1 = 7.818132904e-7   k2 = 5.099082976e-02 wk2 = -3.023925866e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.533532193e+05 wvsat = -5.512476901e-1   ua = -1.513984172e-09 wua = 1.239354524e-15   ub = 2.952053795e-18 wub = -1.345493439e-24   uc = 7.260003938e-11 wuc = -1.078016999e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.171789723e-02 wu0 = 4.058406654e-9   a0 = 2.279338622e+00 wa0 = -1.793266905e-6   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 6.229599982e-01 wags = -2.468558888e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.250892197e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 3.088599517e-8   nfactor = {5.552014819e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.086907266e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.754532663e-05 wcit = -3.767411769e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.300775800e-01 wpclm = 9.912361758e-7   pdiblc1 = 0.39   pdiblc2 = 6.399121367e-03 wpdiblc2 = 9.380855305e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.619336596e-05 walpha0 = 3.793003797e-11   alpha1 = 0.0   beta0 = 1.715745884e+01 wbeta0 = 1.916813899e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.513589544e-01 wkt1 = -1.333663766e-8   kt2 = -3.455418412e-02 wkt2 = -6.781341185e-10   at = -3.097523218e+05 wat = 1.886606792e+0   ute = -1.100168913e+00 wute = -4.829821888e-7   ua1 = 4.193518501e-09 wua1 = -6.332265702e-15   ub1 = -5.060436973e-18 wub1 = 8.924244999e-24   uc1 = 2.967892342e-12 wuc1 = -1.495210383e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.26 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.237426502e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.424717146e-08 wvth0 = 7.320856975e-09 pvth0 = 9.767756566e-14   k1 = -7.952435560e-02 lk1 = 1.277400177e-06 wk1 = 1.933047248e-06 pk1 = -4.549325473e-12   k2 = 1.716357775e-01 lk2 = -4.767520367e-07 wk2 = -7.449097288e-07 pk2 = 1.748692778e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.352633700e+05 lvsat = -1.114022933e+00 wvsat = -1.011954505e+00 pvsat = 1.820572818e-6   ua = -1.746498130e-09 lua = 9.188242437e-16 wua = 2.333584938e-15 pua = -4.324064854e-21   ub = 3.098022211e-18 lub = -5.768226571e-25 wub = -2.157540947e-24 pub = 3.208964075e-30   uc = 3.854774482e-11 luc = 1.345642822e-16 wuc = 3.315515159e-17 puc = -1.736189906e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.944981847e-02 lu0 = 8.962755520e-09 wu0 = 1.268387469e-08 pu0 = -3.408521892e-14   a0 = 2.521425850e+00 la0 = -9.566548864e-07 wa0 = -3.081978358e-06 pa0 = 5.092594606e-12   keta = 1.580486228e-01 lketa = -6.245599525e-07 wketa = 2.633051543e-07 pketa = -1.040501662e-12   a1 = 0.0   a2 = 0.38689047   ags = 3.777367213e-01 lags = 9.690475974e-07 wags = -3.263218267e-06 pags = 1.191974413e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.481449664e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.110927916e-08 wvoff = 1.092036538e-07 pvoff = -3.094875000e-13   nfactor = {-5.219941464e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.256748578e-06 wnfactor = 5.254696946e-06 pnfactor = -1.251813864e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.978765226e-05 lcit = -4.837793699e-11 wcit = -7.443831126e-11 pcit = 1.452808799e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378098707e-01 letab = 2.679639268e-07 wetab = -5.757272712e-11 petab = 2.275098579e-16   dsub = 5.817163284e-01 ldsub = -8.581630639e-08 wdsub = 5.671023179e-07 pdsub = -2.241015394e-12   voffl = 0.0   minv = 0.0   pclm = -1.071292677e-01 lpclm = -9.068473084e-08 wpclm = 9.699129435e-07 ppclm = 8.426291034e-14   pdiblc1 = 0.39   pdiblc2 = 2.893893137e-03 lpdiblc2 = 1.385159287e-08 wpdiblc2 = 7.737990772e-09 ppdiblc2 = -2.687115154e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.520959765e-05 lalpha0 = 3.216796843e-10 walpha0 = -2.000617673e-11 palpha0 = 2.289462500e-16   alpha1 = 0.0   beta0 = 1.332170879e+01 lbeta0 = 1.515771429e-05 wbeta0 = 2.670273988e-06 pbeta0 = -2.977444465e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.220327527e-01 lkt1 = -1.158882044e-07 wkt1 = -1.082617854e-07 pkt1 = 3.751152319e-13   kt2 = -6.815623071e-02 lkt2 = 1.327850395e-07 wkt2 = 1.045262822e-07 pkt2 = -4.157357659e-13   at = -6.916769417e+05 lat = 1.509249611e+00 wat = 3.841638371e+00 pat = -7.725688518e-6   ute = -9.361382218e-01 lute = -6.481992605e-07 wute = -1.124149725e-06 pute = 2.533698545e-12   ua1 = 5.129144791e-09 lua1 = -3.697309735e-15 wua1 = -9.563103032e-15 pua1 = 1.276728372e-20   ub1 = -6.639192552e-18 lub1 = 6.238760526e-24 wub1 = 1.486975038e-23 pub1 = -2.349482390e-29   uc1 = 2.381160033e-11 luc1 = -8.236797663e-17 wuc1 = -1.925866146e-16 puc1 = 1.701820227e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.27 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.073713932e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.770452900e-08 wvth0 = 8.057799350e-08 pvth0 = -4.529802141e-14   k1 = 7.107031071e-01 lk1 = -2.648828104e-07 wk1 = -7.918807436e-07 pk1 = 7.689028631e-13   k2 = -1.189729771e-01 lk2 = 9.042761654e-08 wk2 = 2.998843880e-07 pk2 = -2.904266754e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.136687958e+04 lvsat = 6.047977934e-03 wvsat = -1.842486279e-01 pvsat = 2.051433958e-7   ua = -9.699709012e-10 lua = -5.967200655e-16 wua = -7.655214051e-17 pua = 3.797876312e-22   ub = 2.762828214e-18 lub = 7.737379057e-26 wub = -6.900373675e-25 pub = 3.448446769e-31   uc = 1.335007973e-10 luc = -5.075511562e-17 wuc = -8.991465507e-17 puc = 6.657573571e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.816167661e-02 lu0 = -8.040134451e-09 wu0 = -7.510344800e-09 pu0 = 5.327738295e-15   a0 = 1.946997424e+00 la0 = 1.644542005e-07 wa0 = 6.079738586e-07 pa0 = -2.109066685e-12   keta = -1.786231207e-01 lketa = 3.252060604e-08 wketa = -4.094385561e-07 pketa = 2.724888741e-13   a1 = 0.0   a2 = 0.38689047   ags = -1.866657576e-01 lags = 2.070589093e-06 wags = 5.206707682e-06 pags = -4.610967998e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.883957187e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.463676288e-08 wvoff = -9.243037975e-08 pvoff = 8.404063509e-14   nfactor = {1.843830718e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.606199796e-07 wnfactor = -3.133201742e-06 pnfactor = 3.852481291e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.163487279e-04 leta0 = -3.190773040e-11 weta0 = 4.861838936e-11 peta0 = -9.488826742e-17   etab = -5.404702030e-04 letab = 5.592430080e-11 wetab = 8.954550587e-11 petab = -5.962006183e-17   dsub = -2.105686038e-01 ldsub = 1.460482234e-06 wdsub = 4.055997035e-07 pdsub = -1.925811549e-12   voffl = 0.0   minv = 0.0   pclm = -8.232740390e-01 lpclm = 1.307011439e-06 wpclm = 3.292013213e-06 ppclm = -4.447768575e-12   pdiblc1 = 0.39   pdiblc2 = 9.778393952e-03 lpdiblc2 = 4.151470518e-10 wpdiblc2 = -2.038114916e-08 ppdiblc2 = 2.800883327e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.390081162e-04 lalpha0 = -5.737405676e-11 walpha0 = 2.797917887e-10 palpha0 = -3.561679401e-16   alpha1 = 0.0   beta0 = 2.034063118e+01 lbeta0 = 1.458918552e-06 wbeta0 = 5.267107457e-06 pbeta0 = -8.045671362e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.986870767e-01 lkt1 = 3.371765636e-08 wkt1 = 1.693428040e-07 pkt1 = -1.666842574e-13   kt2 = 5.475960451e-02 lkt2 = -1.071091815e-07 wkt2 = -3.170148204e-07 pkt2 = 4.069838962e-13   at = 9.396629926e+04 lat = -2.408637446e-02 wat = -2.522052616e-01 pat = 2.642456308e-7   ute = -1.263602351e+00 lute = -9.089156403e-09 wute = -1.371606350e-07 pute = 6.073968740e-13   ua1 = 4.993351616e-09 lua1 = -3.432282873e-15 wua1 = -9.648767402e-15 pua1 = 1.293447445e-20   ub1 = -5.956811982e-18 lub1 = 4.906961780e-24 wub1 = 1.198231333e-23 pub1 = -1.785942744e-29   uc1 = -9.492617849e-11 luc1 = 1.493719526e-16 wuc1 = 2.225837674e-16 puc1 = -6.401039361e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.28 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.287844838e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.674202310e-09 wvth0 = 5.617671065e-08 pvth0 = -2.207544253e-14   k1 = 4.040518093e-01 lk1 = 2.695569643e-08 wk1 = 1.195818834e-07 pk1 = -9.853156172e-14   k2 = -3.512017179e-03 lk2 = -1.945600168e-08 wk2 = -6.467781921e-08 pk2 = 5.652535441e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -6.391885541e+04 lvsat = 1.252817855e-01 wvsat = 2.063230085e-01 pvsat = -1.665616776e-7   ua = -1.085419338e-09 lua = -4.868483658e-16 wua = -1.846577356e-15 pua = 2.064311778e-21   ub = 2.595657059e-18 lub = 2.364697428e-25 wub = 1.744121879e-24 pub = -1.971732508e-30   uc = 9.196755887e-11 luc = -1.122814027e-17 wuc = 1.287807784e-17 puc = -3.125159423e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.620826194e-02 lu0 = -6.181079478e-09 wu0 = -1.885336521e-08 pu0 = 1.612283411e-14   a0 = 2.949866282e+00 la0 = -7.899710770e-07 wa0 = -4.703423173e-06 pa0 = 2.945763313e-12   keta = -2.914478577e-01 lketa = 1.398953441e-07 wketa = -1.519603025e-07 pketa = 2.744810752e-14   a1 = 0.0   a2 = 0.38689047   ags = 4.769755569e+00 lags = -2.646412301e-06 wags = -4.458627437e-06 pags = 4.587483109e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.103737273e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.142814852e-09 wvoff = -3.065802576e-08 pvoff = 2.525219466e-14   nfactor = {7.713319884e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.600716985e-07 wnfactor = 1.117977876e-06 pnfactor = -1.933450955e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 9.326303828e-04 leta0 = -4.280808113e-10 weta0 = -1.653056211e-10 peta0 = 1.087021437e-16   etab = -9.093683501e-04 letab = 4.070028229e-10 wetab = 2.982940965e-10 petab = -2.582850518e-16   dsub = 1.616780294e+00 ldsub = -2.785965748e-07 wdsub = -3.079608679e-06 pdsub = 1.391043842e-12   voffl = 0.0   minv = 0.0   pclm = 5.761006626e-01 lpclm = -2.476646814e-08 wpclm = -2.013392959e-06 ppclm = 6.013599523e-13   pdiblc1 = 0.39   pdiblc2 = 1.190975726e-02 lpdiblc2 = -1.613260753e-09 wpdiblc2 = 1.023099817e-08 ppdiblc2 = -1.124594288e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.813049822e-05 lalpha0 = 4.814761789e-11 walpha0 = -1.117477032e-10 palpha0 = 1.645823658e-17   alpha1 = 0.0   beta0 = 1.974222689e+01 lbeta0 = 2.028416919e-06 wbeta0 = -4.743956813e-06 pbeta0 = 1.481808448e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.513901226e-01 lkt1 = -1.129461831e-08 wkt1 = -5.991654380e-08 pkt1 = 5.150071766e-14   kt2 = -6.593508084e-02 lkt2 = 7.755347059e-09 wkt2 = 1.458791327e-07 pkt2 = -3.354996437e-14   at = 1.147141437e+05 lat = -4.383199430e-02 wat = -9.855518311e-02 pat = 1.180176194e-7   ute = -2.158126929e+00 lute = 8.422254121e-07 wute = 4.341509852e-06 pute = -3.654931435e-12   ua1 = -2.408113313e-09 lua1 = 3.611654292e-15 wua1 = 2.186222732e-14 pua1 = -1.705438168e-20   ub1 = 4.175098949e-18 lub1 = -4.735527192e-24 wub1 = -2.984804818e-23 pub1 = 2.195031846e-29   uc1 = 1.771225772e-10 luc1 = -1.095354879e-16 wuc1 = -1.033904331e-15 puc1 = 5.556895045e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.29 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.944466127e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.233345763e-08 wvth0 = 9.227639144e-10 pvth0 = 2.882488943e-15   k1 = 3.393828136e-01 lk1 = 5.616635844e-08 wk1 = -1.110996379e-07 pk1 = 5.666128041e-15   k2 = -1.674027854e-02 lk2 = -1.348086216e-08 wk2 = 7.487639978e-08 pk2 = -6.510588539e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.684478581e+05 lvsat = -2.484659718e-02 wvsat = -3.127663460e-01 pvsat = 6.790838833e-8   ua = -3.032405924e-09 lua = 3.925957402e-16 wua = 7.526049717e-15 pua = -2.169257007e-21   ub = 3.807659289e-18 lub = -3.109856044e-25 wub = -6.489405188e-24 pub = 1.747310501e-30   uc = 5.352129683e-11 luc = 6.137844064e-18 wuc = -1.343320403e-17 puc = -1.936691977e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.253839190e-02 lu0 = 4.510482471e-09 wu0 = 6.238906851e-08 pu0 = -2.057396699e-14   a0 = 1.061757793e+00 la0 = 6.287808685e-08 wa0 = 2.991768010e-06 pa0 = -5.301160684e-13   keta = 6.416271625e-02 lketa = -2.073217413e-08 wketa = -1.778311095e-07 pketa = 3.913382171e-14   a1 = 0.0   a2 = 0.38689047   ags = -1.967750237e+00 lags = 3.968853840e-07 wags = 1.029417355e-05 pags = -2.076283335e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.243600741e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.174748096e-09 wvoff = 3.865650442e-08 pvoff = -6.056832054e-15   nfactor = {2.358017877e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.662638404e-08 wnfactor = 5.789960921e-07 pnfactor = 5.011028150e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.706794045e-03 leta0 = -1.229461586e-09 weta0 = -2.795736408e-08 peta0 = 1.266223599e-14   etab = 9.118507360e-02 letab = -4.119159613e-08 wetab = -2.292852444e-07 petab = 1.034434514e-13   dsub = 1.441167857e+00 ldsub = -1.992733153e-07 wdsub = 4.579122716e-07 pdsub = -2.068366835e-13   voffl = 0.0   minv = 0.0   pclm = 5.884537207e-01 lpclm = -3.034628268e-08 wpclm = -1.048961173e-06 ppclm = 1.657309365e-13   pdiblc1 = 0.39   pdiblc2 = 5.686669736e-03 lpdiblc2 = 1.197676767e-09 wpdiblc2 = 7.286068271e-10 ppdiblc2 = 3.167588371e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.042076695e-03 lalpha0 = 5.315548560e-10 walpha0 = -1.144884246e-09 palpha0 = 4.831208475e-16   alpha1 = 0.0   beta0 = 1.914616876e+01 lbeta0 = 2.297653399e-06 wbeta0 = -2.479489381e-06 pbeta0 = 4.589598311e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.320547566e-01 lkt1 = 2.514119353e-08 wkt1 = 2.518481117e-07 pkt1 = -8.932181842e-14   kt2 = -5.821091455e-02 lkt2 = 4.266379767e-09 wkt2 = 8.458805447e-08 pkt2 = -5.865090813e-15   at = 2.092526313e+03 lat = 7.038627176e-03 wat = 2.470005417e-01 pat = -3.806817370e-8   ute = -8.907282010e-01 lute = 2.697477434e-07 wute = -1.594730959e-06 pute = -9.735611416e-13   ua1 = 4.976047728e-09 lua1 = 2.762656707e-16 wua1 = -1.337449054e-14 pua1 = -1.138132405e-21   ub1 = -6.530591402e-18 lub1 = 1.001796105e-25 wub1 = 1.910189420e-23 pub1 = -1.601257658e-31   uc1 = -1.548287735e-10 luc1 = 4.040527742e-17 wuc1 = 5.380066200e-16 puc1 = -1.543348124e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.30 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.243303493e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.853035788e-08 wvth0 = -1.913091876e-07 pvth0 = 4.165471240e-14   k1 = 4.246445314e-01 lk1 = 3.896949628e-08 wk1 = -8.012176134e-08 pk1 = -5.819547735e-16   k2 = -6.255996722e-02 lk2 = -4.239260056e-09 wk2 = 5.689326898e-08 pk2 = -2.883480971e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.031315822e+05 lvsat = 8.496869102e-03 wvsat = 1.649119128e-01 pvsat = -2.843692809e-8   ua = 1.886895471e-09 lua = -5.996027546e-16 wua = -1.179086314e-14 pua = 1.726867732e-21   ub = 9.588450248e-19 lub = 2.636059886e-25 wub = 7.975708443e-24 pub = -1.170230593e-30   uc = 1.839357345e-10 luc = -2.016609594e-17 wuc = -3.616169289e-16 puc = 5.085999661e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.760132598e-02 lu0 = -8.612386020e-09 wu0 = -1.332387497e-07 pu0 = 1.888318580e-14   a0 = 3.957561783e+00 la0 = -5.211910991e-07 wa0 = 1.047265436e-06 pa0 = -1.379196216e-13   keta = -2.796445986e-02 lketa = -2.150583345e-09 wketa = 4.234236939e-07 pketa = -8.213626586e-14   a1 = 0.0   a2 = 0.38689047   ags = -2.385479756e+00 lags = 4.811393395e-07 wags = 7.144549818e-07 pags = -1.441019976e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.632928372e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.002729173e-08 wvoff = 5.459487905e-08 pvoff = -9.271522523e-15   nfactor = {-2.041526498e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.601506004e-07 wnfactor = 4.997142952e-06 pnfactor = -8.410078495e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.318630225e-06 lcit = -8.710461233e-13 wcit = -1.296901931e-11 pcit = 2.615786350e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.115436827e-01 leta0 = 4.198378826e-08 weta0 = 2.532998239e-07 peta0 = -4.406593253e-14   etab = -2.875635259e-01 letab = 3.520010264e-08 wetab = 7.862308516e-07 petab = -1.013810676e-13   dsub = 7.570655415e-01 ldsub = -6.129329874e-08 wdsub = -1.882797735e-06 pdsub = 2.652728212e-13   voffl = 0.0   minv = 0.0   pclm = 1.214130247e+00 lpclm = -1.565421097e-07 wpclm = -1.704698865e-06 ppclm = 2.979899503e-13   pdiblc1 = -7.660564720e-01 lpdiblc1 = 2.331708101e-07 wpdiblc1 = 4.209812575e-08 ppdiblc1 = -8.490981473e-15   pdiblc2 = 2.060437795e-02 lpdiblc2 = -1.811150390e-09 wpdiblc2 = 1.649015291e-08 ppdiblc2 = -1.143666647e-17   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.258172791e-04 lalpha0 = 4.879364131e-10 walpha0 = 1.679214769e-08 palpha0 = -3.134688809e-15   alpha1 = 0.0   beta0 = 2.587452690e+01 lbeta0 = 9.405772028e-07 wbeta0 = 2.408760758e-05 pbeta0 = -4.899490791e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 2.081365242e-03 lkt1 = -4.225239156e-08 wkt1 = -6.423618763e-07 pkt1 = 9.103586513e-14   kt2 = -2.149268130e-02 lkt2 = -3.139504289e-09 wkt2 = 2.720018392e-08 pkt2 = 5.709755737e-15   at = -8.540323236e+04 lat = 2.468608422e-02 wat = 3.464085893e-01 pat = -5.811827985e-8   ute = 3.893612047e+00 lute = -6.952297630e-07 wute = -1.659212219e-05 pute = 2.051337682e-12   ua1 = 1.685366291e-08 lua1 = -2.119389924e-15 wua1 = -5.035838573e-14 pua1 = 6.321334336e-21   ub1 = -1.593008240e-17 lub1 = 1.996009946e-24 wub1 = 4.707606220e-23 pub1 = -5.802375580e-30   uc1 = 1.141303070e-10 luc1 = -1.384242432e-17 wuc1 = -5.698571879e-16 puc1 = 6.911577833e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.31 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.524259436e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.617092834e-09 wvth0 = 5.007585555e-07 pvth0 = -4.948714902e-14   k1 = 6.607947852e-01 lk1 = 7.869688600e-09 wk1 = 5.445537152e-07 pk1 = -8.284859165e-14   k2 = -1.514686236e-01 lk2 = 7.469565447e-09 wk2 = -8.564086017e-08 pk2 = 1.588755117e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.429229479e+05 lvsat = -9.912954803e-03 wvsat = -2.277930602e-01 pvsat = 2.328035334e-8   ua = -2.997406310e-09 lua = 4.363536840e-17 wua = 3.879105399e-15 pua = -3.367887753e-22   ub = 1.808014123e-18 lub = 1.517746642e-25 wub = 3.575724488e-24 pub = -5.907747057e-31   uc = 1.019392468e-10 luc = -9.367568493e-18 wuc = -7.510581935e-17 puc = 1.312791604e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -5.607839414e-03 lu0 = 2.345845017e-09 wu0 = 9.509671087e-08 pu0 = -1.118745268e-14   a0 = 0.0   keta = -2.346717703e-01 lketa = 2.507173590e-08 wketa = 1.032478670e-06 pketa = -1.623457610e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.300217953e+00 lags = -4.248620411e-09 wags = -1.554677722e-06 pags = 1.547314339e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {1.423370787e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.022264004e-08 wvoff = -8.073134982e-07 pvoff = 1.042375012e-13   nfactor = {5.603822195e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.047306468e-07 wnfactor = -1.402417827e-05 pnfactor = 1.664005049e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.050059587e-05 lcit = -2.343655089e-12 wcit = -9.744793490e-11 pcit = 1.374123714e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.541029829e-01 leta0 = -3.250904936e-08 weta0 = -8.120423143e-07 peta0 = 9.623430036e-14   etab = 1.170738274e-02 letab = -4.212379674e-09 wetab = -2.304324678e-07 petab = 3.250840824e-14   dsub = 3.989249251e-01 ldsub = -1.412797025e-08 wdsub = 5.772591178e-07 pdsub = -5.870436599e-14   voffl = 0.0   minv = 0.0   pclm = -1.312125510e+00 lpclm = 1.761531423e-07 wpclm = 5.015327850e-06 ppclm = -5.870039679e-13   pdiblc1 = 1.977907512e+00 lpdiblc1 = -1.281955268e-07 wpdiblc1 = -2.975864244e-06 ppdiblc1 = 3.889595729e-13   pdiblc2 = 3.499971289e-02 lpdiblc2 = -3.706944026e-09 wpdiblc2 = -2.157912304e-09 ppdiblc2 = 2.444420282e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.850201331e-03 lalpha0 = -7.863468578e-10 walpha0 = -2.279940534e-08 palpha0 = 2.079320768e-15   alpha1 = 0.0   beta0 = 3.989051912e+01 lbeta0 = -9.052588925e-07 wbeta0 = -2.677712182e-05 pbeta0 = 1.799139747e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -8.690562389e-01 lkt1 = 7.247207522e-08 wkt1 = 2.243962952e-06 pkt1 = -2.890786832e-13   kt2 = -1.569903007e-01 lkt2 = 1.470485470e-08 wkt2 = 3.021690937e-07 pkt2 = -3.050227483e-14   at = 2.600051028e+05 lat = -2.080246648e-02 wat = -7.386820704e-01 pat = 8.478273458e-8   ute = -2.478690182e+00 lute = 1.439705791e-07 wute = 1.653423468e-06 pute = -3.515094530e-13   ua1 = -3.211823563e-10 lua1 = 1.424513236e-16 wua1 = -9.211904921e-16 pua1 = -1.892970907e-22   ub1 = 1.472021668e-19 lub1 = -1.212880440e-25 wub1 = 3.410083946e-24 pub1 = -5.178457444e-32   uc1 = 5.860431172e-11 luc1 = -6.529928377e-18 wuc1 = 1.443369310e-16 puc1 = -2.494001616e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.32 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.43080609+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.50407   k2 = -0.049704661   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169790.0   ua = -1.1012842e-9   ub = 2.50401e-18   uc = 6.9010287e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03306933   a0 = 1.6821881   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.540758   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.25013304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0067115   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.8823913e-5   alpha1 = 0.0   beta0 = 17.79575   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.2558   kt2 = -0.03478   at = 318480.0   ute = -1.261   ua1 = 2.0849e-9   ub1 = -2.0887e-18   uc1 = -4.6822e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.33 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.43080609+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.50407   k2 = -0.049704661   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169790.0   ua = -1.1012842e-9   ub = 2.50401e-18   uc = 6.9010287e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03306933   a0 = 1.6821881   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.540758   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.25013304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0067115   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.8823913e-5   alpha1 = 0.0   beta0 = 17.79575   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.2558   kt2 = -0.03478   at = 318480.0   ute = -1.261   ua1 = 2.0849e-9   ub1 = -2.0887e-18   uc1 = -4.6822e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.34 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.261804655e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.827905718e-8   k1 = 5.641724475e-01 lk1 = -2.375065414e-7   k2 = -7.641610622e-02 lk2 = 1.055554845e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.982866713e+05 lvsat = -5.077796533e-1   ua = -9.694239190e-10 lua = -5.210716130e-16   ub = 2.379569927e-18 lub = 4.917492151e-25   uc = 4.958827428e-11 luc = 7.674987057e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.367349670e-02 lu0 = -2.387482544e-9   a0 = 1.495139700e+00 la0 = 7.391582251e-7   keta = 2.457281590e-01 lketa = -9.710427372e-7   a1 = 0.0   a2 = 0.38689047   ags = -7.089015742e-01 lags = 4.938273491e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.117805977e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.194878866e-8   nfactor = {1.227798379e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.825976766e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378290421e-01 letab = 2.680396867e-7   dsub = 7.705590737e-01 ldsub = -8.320652388e-7   voffl = 0.0   minv = 0.0   pclm = 2.158477634e-01 lpclm = -6.262552739e-8   pdiblc1 = 0.39   pdiblc2 = 5.470612319e-03 lpdiblc2 = 4.903609645e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.187157242e-05 lalpha0 = 3.979178463e-10   alpha1 = 0.0   beta0 = 1.421089907e+01 lbeta0 = 1.416623750e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.580834831e-01 lkt1 = 9.023628946e-9   kt2 = -3.334940756e-02 lkt2 = -5.653264972e-9   at = 5.875728757e+05 lat = -1.063372971e+0   ute = -1.310475468e+00 lute = 1.955119605e-7   ua1 = 1.944670714e-09 lua1 = 5.541433674e-16   ub1 = -1.687626677e-18 lub1 = -1.584919443e-24   uc1 = -4.031895226e-11 luc1 = -2.569806124e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.35 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.342035344e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.620473702e-9   k1 = 4.470100682e-01 lk1 = -8.841311456e-9   k2 = -1.911270615e-02 lk2 = -6.283274872e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.284237000e+01 lvsat = 7.435988715e-2   ua = -9.954624500e-10 lua = -4.702523424e-16   ub = 2.533048601e-18 lub = 1.922056532e-25   uc = 1.035595861e-10 luc = -2.858566876e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.566076260e-02 lu0 = -6.266019456e-9   a0 = 2.149450225e+00 la0 = -5.378563531e-7   keta = -3.149644802e-01 lketa = 1.232582832e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.547146540e+00 lags = 5.351556668e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.196185091e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.348423824e-9   nfactor = {8.004873916e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.222404856e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.325384520e-04 leta0 = -6.350513417e-11   etab = -5.106519169e-04 letab = 3.607106480e-11   dsub = -7.550556647e-02 ldsub = 8.191948891e-7   voffl = 0.0   minv = 0.0   pclm = 2.729528554e-01 lpclm = -1.740772499e-7   pdiblc1 = 0.39   pdiblc2 = 2.991554895e-03 lpdiblc2 = 9.741973625e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.321776340e-04 lalpha0 = -1.759765196e-10   alpha1 = 0.0   beta0 = 2.209455635e+01 lbeta0 = -1.220257004e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.422966176e-01 lkt1 = -2.178751752e-8   kt2 = -5.080503011e-02 lkt2 = 2.841478627e-8   at = 9.982981830e+03 lat = 6.390633654e-2   ute = -1.309276280e+00 lute = 1.931715108e-7   ua1 = 1.780351655e-09 lua1 = 8.748440537e-16   ub1 = -1.966750800e-18 lub1 = -1.040154289e-24   uc1 = -2.080669709e-11 luc1 = -6.378003209e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.36 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.474910980e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.002523411e-8   k1 = 4.438720859e-01 lk1 = -5.854909391e-9   k2 = -2.504946564e-02 lk2 = -6.332905569e-10   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.785859965e+03 lvsat = 6.981743017e-02 pvsat = 6.776263578e-21   ua = -1.700322021e-09 lua = 2.005589875e-16   ub = 3.176442490e-18 lub = -4.201090932e-25   uc = 9.625590596e-11 luc = -2.163479294e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.993016867e-02 lu0 = -8.122418646e-10   a0 = 1.383645661e+00 la0 = 1.909560213e-7   keta = -3.420500150e-01 lketa = 1.490354513e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.285050924e+00 lags = -1.118799246e-06 wags = -4.336808690e-19   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.205827241e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.266062371e-9   nfactor = {1.143614035e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.956885749e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.775841959e-04 leta0 = -3.918834434e-10   etab = -8.100376397e-04 letab = 3.209949603e-10   dsub = 5.912832380e-01 ldsub = 1.846153178e-7   voffl = 0.0   minv = 0.0   pclm = -9.435093290e-02 lpclm = 1.754839289e-07 ppclm = -1.292469707e-26   pdiblc1 = 0.39   pdiblc2 = 1.531663768e-02 lpdiblc2 = -1.987746037e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -9.081028498e-06 lalpha0 = 5.362814315e-11   alpha1 = 0.0   beta0 = 1.816250874e+01 lbeta0 = 2.521853053e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.713420859e-01 lkt1 = 5.854909391e-9   kt2 = -1.735792814e-02 lkt2 = -3.416653439e-9   at = 8.189567208e+04 lat = -4.532611205e-3   ute = -7.124219600e-01 lute = -3.748517613e-7   ua1 = 4.871918696e-09 lua1 = -2.067384841e-15   ub1 = -5.764178643e-18 lub1 = 2.573838802e-24   uc1 = -1.671633234e-10 luc1 = 7.550683735e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.37 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.947538893e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.137360064e-8   k1 = 3.023870900e-01 lk1 = 5.805315583e-8   k2 = 8.193255407e-03 lk2 = -1.564886144e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.642979480e+05 lvsat = -2.233382459e-3   ua = -5.262622437e-10 lua = -3.297579438e-16   ub = 1.646713984e-18 lub = 2.708616242e-25   uc = 4.904809500e-11 luc = -3.112607667e-19   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.331369576e-02 lu0 = -2.340564133e-9   a0 = 2.058004266e+00 la0 = -1.136483891e-7   keta = 4.945686336e-03 lketa = -7.700772046e-9   a1 = 0.0   a2 = 0.38689047   ags = 1.460167325e+00 lags = -2.945084486e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.114876168e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.578478699e-10   nfactor = {2.550821201e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.993986587e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -6.602893771e-03 leta0 = 2.987011052e-09 weta0 = -1.257314531e-22 peta0 = -1.494891415e-28   etab = 1.483402786e-02 letab = -6.745351206e-09 wetab = -2.646977960e-22 petab = 1.262177448e-28   dsub = 1.593650765e+00 ldsub = -2.681490824e-7   voffl = 0.0   minv = 0.0   pclm = 2.391539534e-01 lpclm = 2.484143925e-8   pdiblc1 = 0.39   pdiblc2 = 5.929292820e-03 lpdiblc2 = 2.252470700e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.423318452e-03 lalpha0 = 6.924321162e-10 walpha0 = 7.940933881e-23 palpha0 = 3.786532345e-29   alpha1 = 0.0   beta0 = 1.832050896e+01 lbeta0 = 2.450485140e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.481903686e-01 lkt1 = -4.602605555e-9   kt2 = -3.004343944e-02 lkt2 = 2.313328588e-9   at = 8.434269338e+04 lat = -5.637918491e-3   ute = -1.421767068e+00 lute = -5.444412272e-8   ua1 = 5.223972481e-10 lua1 = -1.027277508e-16   ub1 = -1.697389995e-19 lub1 = 4.685838739e-26 pub1 = 2.802596929e-45   uc1 = 2.432522378e-11 luc1 = -1.098758196e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.38 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.606251747e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.465950954e-8   k1 = 3.979643136e-01 lk1 = 3.877570772e-8   k2 = -4.361474206e-02 lk2 = -5.199447390e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.580465726e+05 lvsat = -9.725112878e-4   ua = -2.039413583e-09 lua = -2.456288450e-17   ub = 3.614723216e-18 lub = -1.260759979e-25   uc = 6.351878069e-11 luc = -3.229925718e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.323336894e-02 lu0 = -2.324362616e-9   a0 = 4.306296877e+00 la0 = -5.671177672e-7   keta = 1.130338931e-01 lketa = -2.950162291e-8   a1 = 0.0   a2 = 0.38689047   ags = -2.147569179e+00 lags = 4.331539655e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.451129664e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.939912769e-9   nfactor = {1.459875453e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.800984368e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.271958805e-01 leta0 = 2.731001350e-08 weta0 = 6.776263578e-21 peta0 = -8.077935669e-28   etab = -2.575187780e-02 letab = 1.440623036e-9   dsub = 1.301016200e-01 ldsub = 2.704146245e-8   voffl = 0.0   minv = 0.0   pclm = 6.464725184e-01 lpclm = -5.731267872e-8   pdiblc1 = -7.520379688e-01 lpdiblc1 = 2.303433481e-7   pdiblc2 = 2.609553121e-02 lpdiblc2 = -1.814958753e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.765899011e-03 lalpha0 = -5.559021000e-10   alpha1 = 0.0   beta0 = 3.389560141e+01 lbeta0 = -6.909331302e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.118225043e-01 lkt1 = -1.193782195e-8   kt2 = -1.243513164e-02 lkt2 = -1.238179053e-9   at = 2.994940671e+04 lat = 5.332935463e-3   ute = -1.631496571e+00 lute = -1.214273053e-8   ua1 = 8.452706293e-11 lua1 = -1.441152383e-17 wua1 = 6.310887242e-30 pua1 = 7.523163845e-37   ub1 = -2.539468139e-19 lub1 = 6.384268250e-26 wub1 = 2.350988702e-38 pub1 = 2.802596929e-45   uc1 = -7.562979876e-11 luc1 = 9.172846315e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.39 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.803347206e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.666638331e-07 wvth0 = 6.374023555e-06 pvth0 = -8.394270320e-13   k1 = 8.421289383e-01 lk1 = -1.971855253e-8   k2 = 7.148822975e-01 lk2 = -1.050897150e-07 wk2 = -2.687327330e-06 pk2 = 3.539075728e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.355540881e+06 lvsat = -2.903715243e-01 wvsat = -6.572069220e+00 pvsat = 8.655086559e-7   ua = 3.188609819e-08 lua = -4.492383157e-15 wua = -1.008774539e-13 pua = 1.328505630e-20   ub = -3.531121363e-17 lub = 5.000275255e-24 wub = 1.150462502e-22 pub = -1.515101592e-29   uc = 7.692931709e-11 luc = -4.996026308e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.548105320e-01 lu0 = -1.833546710e-08 wu0 = -3.866460751e-07 pu0 = 5.091935486e-14   a0 = 0.0   keta = 1.091393912e-01 lketa = -2.898873649e-8   a1 = 0.0   a2 = 0.38689047   ags = 7.825166500e-01 lags = 4.727631228e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.264950042e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.488020234e-9   nfactor = {-4.634609714e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.475905997e-06 wnfactor = 1.419835075e-04 pnfactor = -1.869851802e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.194916667e-05 lcit = 2.232120504e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.369622363e-02 leta0 = -4.634221449e-10   etab = -6.502568369e-02 letab = 6.612786903e-9   dsub = 5.911498431e-01 ldsub = -3.367628329e-8   voffl = 0.0   minv = 0.0   pclm = 3.579580883e-01 lpclm = -1.931677084e-8   pdiblc1 = 9.869569272e-01 lpdiblc1 = 1.326415288e-9   pdiblc2 = 3.428113695e-02 lpdiblc2 = -2.892962101e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.258092888e-03 lalpha0 = -9.394157264e-11   alpha1 = 0.0   beta0 = 3.097384741e+01 lbeta0 = -3.061527377e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.218257817e-01 lkt1 = -2.378994033e-8   kt2 = -5.636923217e-02 lkt2 = 4.547722315e-9   at = 1.402700383e+04 lat = 7.429836310e-3   ute = -1.928106950e+00 lute = 2.691937328e-8   ua1 = -6.279350110e-10 lua1 = 7.941616899e-17 wua1 = 2.524354897e-29 pua1 = -4.513898307e-36   ub1 = 1.282746131e-18 lub1 = -1.385320949e-25 pub1 = 1.121038771e-44   uc1 = 1.066679176e-10 luc1 = -1.483485144e-17 wuc1 = -3.155443621e-30 puc1 = 3.761581923e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.40 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.394666025e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.592126040e-8   k1 = 4.685438240e-01 wk1 = 1.063312658e-7   k2 = -4.055360124e-02 wk2 = -2.738948791e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.323530293e+05 wvsat = 1.120503507e-1   ua = -1.248192666e-09 wua = 4.397029155e-16   ub = 2.639359984e-18 wub = -4.051079161e-25   uc = 1.257982525e-10 wuc = -1.699686524e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.300383964e-02 wu0 = 1.960152591e-10   a0 = 1.389379751e+00 wa0 = 8.763871013e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.793689532e-01 wags = -1.155641273e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.203665724e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.664807392e-8   nfactor = {8.901286633e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.077507500e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.085333333e-06 wcit = 1.821364608e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 5.667743627e-03 wpdiblc2 = 3.124004576e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.528100272e-05 walpha0 = 1.060407217e-11   alpha1 = 0.0   beta0 = 1.779865514e+01 wbeta0 = -8.695194639e-9   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.535727680e-01 wkt1 = -6.666194465e-9   kt2 = -3.285216640e-02 wkt2 = -5.770083078e-9   at = 6.352216000e+05 wat = -9.480202785e-1   ute = -1.358608747e+00 wute = 2.921468831e-7   ua1 = 2.232530187e-09 wua1 = -4.418630539e-16   ub1 = -2.846567413e-18 wub1 = 2.268327483e-24   uc1 = -1.809914293e-10 wuc1 = 4.015744688e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.41 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.394666025e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.592126040e-8   k1 = 4.685438240e-01 wk1 = 1.063312658e-7   k2 = -4.055360124e-02 wk2 = -2.738948791e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.323530293e+05 wvsat = 1.120503507e-1   ua = -1.248192666e-09 wua = 4.397029155e-16   ub = 2.639359984e-18 wub = -4.051079161e-25   uc = 1.257982525e-10 wuc = -1.699686524e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.300383964e-02 wu0 = 1.960152591e-10   a0 = 1.389379751e+00 wa0 = 8.763871013e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.793689532e-01 wags = -1.155641273e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.203665724e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.664807392e-8   nfactor = {8.901286633e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.077507500e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.085333333e-06 wcit = 1.821364608e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 5.667743627e-03 wpdiblc2 = 3.124004576e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.528100272e-05 walpha0 = 1.060407217e-11   alpha1 = 0.0   beta0 = 1.779865514e+01 wbeta0 = -8.695194639e-9   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.535727680e-01 wkt1 = -6.666194465e-9   kt2 = -3.285216640e-02 wkt2 = -5.770083078e-9   at = 6.352216000e+05 wat = -9.480202785e-1   ute = -1.358608747e+00 wute = 2.921468831e-7   ua1 = 2.232530187e-09 wua1 = -4.418630539e-16   ub1 = -2.846567413e-18 wub1 = 2.268327483e-24   uc1 = -1.809914293e-10 wuc1 = 4.015744688e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.42 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.380677508e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.527835543e-09 wvth0 = -3.557912023e-08 pvth0 = 3.816491641e-14   k1 = 5.123276656e-01 lk1 = -1.730203880e-07 wk1 = 1.551735061e-07 pk1 = -1.930096366e-13   k2 = -6.433215472e-02 lk2 = 9.396559092e-08 wk2 = -3.616775019e-08 pk2 = 3.468901514e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.297624000e+05 lvsat = -3.849321231e-01 wvsat = 2.050958848e-01 pvsat = -3.676875719e-7   ua = -1.111959640e-09 lua = -5.383513677e-16 wua = 4.266151147e-16 pua = 5.171899707e-23   ub = 2.585443842e-18 lub = 2.130601474e-25 wub = -6.161888641e-25 pub = 8.341275269e-31   uc = 1.173167130e-10 luc = 3.351645723e-17 wuc = -2.027139264e-16 puc = 1.293993355e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.461276453e-02 lu0 = -6.357980427e-09 wu0 = -2.811266169e-09 pu0 = 1.188385898e-14   a0 = 9.075354980e-01 la0 = 1.904101525e-06 wa0 = 1.758722882e-06 pa0 = -3.486721894e-12   keta = 3.295540109e-01 lketa = -1.302296937e-06 wketa = -2.508941279e-07 pketa = 9.914570706e-13   a1 = 0.0   a2 = 0.38689047   ags = -1.032889569e+00 lags = 6.371153942e-06 wags = 9.697090291e-07 pags = -4.288668506e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.217457127e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.449941603e-09 wvoff = 2.982598761e-08 pvoff = -5.207509564e-14   nfactor = {5.387554667e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.388519704e-06 wnfactor = 2.062332999e-06 pnfactor = -3.891730001e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.085333333e-06 wcit = 1.821364608e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378383416e-01 letab = 2.680764353e-07 wetab = 2.783367840e-11 petab = -1.099902077e-16   dsub = 8.394601116e-01 ldsub = -1.104341126e-06 wdsub = -2.062235624e-07 pdsub = 8.149326203e-13   voffl = 0.0   minv = 0.0   pclm = 2.761458436e-01 lpclm = -3.009051495e-07 wpclm = -1.804745660e-07 ppclm = 7.131804403e-13   pdiblc1 = 0.39   pdiblc2 = 7.879773193e-03 lpdiblc2 = -8.741266177e-09 wpdiblc2 = -7.210714862e-09 ppdiblc2 = 4.083965913e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.974723912e-05 lalpha0 = 4.940734781e-10 walpha0 = 8.343298544e-11 palpha0 = -2.877976524e-16   alpha1 = 0.0   beta0 = 1.388635725e+01 lbeta0 = 1.546020802e-05 wbeta0 = 9.713666575e-07 pbeta0 = -3.872905521e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.715691446e-01 lkt1 = 7.111619150e-08 wkt1 = 4.036312420e-08 pkt1 = -1.858455234e-13   kt2 = -3.054150941e-02 lkt2 = -9.131011673e-09 wkt2 = -8.404151493e-09 pkt2 = 1.040903499e-14   at = 1.221060517e+06 lat = -2.315056718e+00 wat = -1.896053849e+00 pat = 3.746339522e-6   ute = -1.395732432e+00 lute = 1.467014805e-07 wute = 2.551775019e-07 pute = 1.460917191e-13   ua1 = 2.019852942e-09 lua1 = 8.404356059e-16 wua1 = -2.250234138e-16 pua1 = -8.568841216e-22   ub1 = -2.466040807e-18 lub1 = -1.503725087e-24 wub1 = 2.329824627e-24 pub1 = -2.430179558e-31   uc1 = -2.528083074e-10 luc1 = 2.837983979e-16 wuc1 = 6.359891395e-16 puc1 = -9.263352821e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.43 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.426655118e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.445591763e-09 wvth0 = -2.532703687e-08 pvth0 = 1.815597658e-14   k1 = 4.331985589e-01 lk1 = -1.858450602e-08 wk1 = 4.133839984e-08 pk1 = 2.916177107e-14   k2 = -1.508700523e-02 lk2 = -2.145921114e-09 wk2 = -1.204908388e-08 pk2 = -1.238326529e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3.987519476e+03 lvsat = 7.127642603e-02 wvsat = 1.197324302e-02 pvsat = 9.228922445e-9   ua = -1.316089196e-09 lua = -1.399527341e-16 wua = 9.596486760e-16 pua = -9.885999395e-22   ub = 2.689080837e-18 lub = 1.079234371e-26 wub = -4.670107216e-25 pub = 5.429772919e-31   uc = 1.589329992e-10 luc = -4.770584037e-17 wuc = -1.657348405e-16 puc = 5.722743845e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.289865482e-02 lu0 = -3.012561075e-09 wu0 = 8.267099076e-09 pu0 = -9.737731072e-15   a0 = 2.053369092e+00 la0 = -3.322161721e-07 wa0 = 2.875746717e-07 pa0 = -6.154892874e-13   keta = -3.981315136e-01 lketa = 1.179232625e-07 wketa = 2.489222575e-07 pketa = 1.596793033e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.909044647e+00 lags = 6.293956425e-07 wags = -1.083175509e-06 pags = -2.820640168e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.205683509e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.152090541e-09 wvoff = 2.842914429e-09 pvoff = 5.876333683e-16   nfactor = {7.266654701e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.021776690e-06 wnfactor = 2.209519637e-07 pnfactor = -2.979158413e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.876714640e-06 lcit = 1.130300994e-11 wcit = 3.554748199e-11 pcit = -3.383036087e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.950913805e-04 leta0 = 9.580128094e-12 weta0 = 1.120805830e-10 peta0 = -2.187471134e-16   etab = -4.910800297e-04 letab = 1.647164557e-11 wetab = -5.857944122e-11 petab = 5.866184575e-17   dsub = -4.594846325e-01 ldsub = 1.430802837e-06 wdsub = 1.149264704e-06 pdsub = -1.830567051e-12   voffl = 0.0   minv = 0.0   pclm = 2.935274057e-01 lpclm = -3.348286573e-07 wpclm = -6.158045196e-08 ppclm = 4.811353923e-13   pdiblc1 = 0.39   pdiblc2 = -4.254498972e-03 lpdiblc2 = 1.494113214e-08 wpdiblc2 = 2.168772907e-08 ppdiblc2 = -1.556128939e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.736846703e-04 lalpha0 = -2.152347622e-10 walpha0 = -1.242322198e-10 palpha0 = 1.175014903e-16   alpha1 = 0.0   beta0 = 2.270945865e+01 lbeta0 = -1.759794880e-06 wbeta0 = -1.840427176e-06 pbeta0 = 1.614858446e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.115508721e-01 lkt1 = -4.602117083e-08 wkt1 = -9.202324618e-08 pkt1 = 7.253229370e-14   kt2 = -5.084813190e-02 lkt2 = 3.050132191e-08 wkt2 = 1.290053792e-10 pkt2 = -6.245084616e-15   at = -3.681351050e+03 lat = 7.526586153e-02 wat = 4.089789488e-02 pat = -3.399951267e-8   ute = -1.508961447e+00 lute = 3.676899843e-07 wute = 5.976656934e-07 pute = -5.223407718e-13   ua1 = 1.397950183e-09 lua1 = 2.054200111e-15 wua1 = 1.144542902e-15 pua1 = -3.529859853e-21   ub1 = -1.859527048e-18 lub1 = -2.687454957e-24 wub1 = -3.209249776e-25 pub1 = 4.930436793e-30   uc1 = -8.216420271e-11 luc1 = -4.924684797e-17 wuc1 = 1.836454686e-16 puc1 = -4.349840140e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.44 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.506172669e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.101323726e-08 wvth0 = -9.356748465e-09 pvth0 = 2.957132953e-15   k1 = 4.442534243e-01 lk1 = -2.910536615e-08 wk1 = -1.141361046e-09 pk1 = 6.958954710e-14   k2 = -2.870753057e-02 lk2 = 1.081666475e-08 wk2 = 1.094873467e-08 pk2 = -3.427017422e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -9.430157648e+03 lvsat = 7.645615757e-02 wvsat = 4.254910936e-02 pvsat = -1.986997667e-8   ua = -2.297171296e-09 lua = 7.937381951e-16 wua = 1.786393753e-15 pua = -1.775409096e-21   ub = 3.720567835e-18 lub = -9.708686754e-25 wub = -1.628588925e-24 pub = 1.648445460e-30   uc = 1.726495124e-10 luc = -6.075977739e-17 wuc = -2.286491198e-16 puc = 1.171026435e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.623042550e-02 lu0 = 3.333559428e-09 wu0 = 1.107347930e-08 pu0 = -1.240854910e-14   a0 = 7.013640118e-01 la0 = 9.544803031e-07 wa0 = 2.042096266e-06 pa0 = -2.285258716e-12   keta = -4.977123622e-01 lketa = 2.126938583e-07 wketa = 4.659036318e-07 pketa = -1.905321587e-13   a1 = 0.0   a2 = 0.38689047   ags = 3.522826175e+00 lags = -9.064321689e-07 wags = -7.116708365e-07 pags = -6.356231563e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.356366405e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.749250639e-08 wvoff = 4.505697394e-08 pvoff = -3.958727600e-14   nfactor = {1.156087498e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.130978933e-07 wnfactor = -3.733357427e-08 pnfactor = -5.210678629e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.921265298e-03 leta0 = -3.251092459e-09 weta0 = -9.109859287e-09 peta0 = 8.557726951e-15   etab = -8.401388808e-04 letab = 3.486692088e-10 wetab = 9.009421854e-11 petab = -8.283013288e-17   dsub = 1.083637219e+00 ldsub = -3.777851349e-08 wdsub = -1.473635158e-06 pdsub = 6.656336328e-13   voffl = 0.0   minv = 0.0   pclm = -3.429381386e-01 lpclm = 2.708924189e-07 wpclm = 7.440314501e-07 ppclm = -2.855614269e-13   pdiblc1 = 0.39   pdiblc2 = 7.997283934e-03 lpdiblc2 = 3.281171604e-09 wpdiblc2 = 2.190711854e-08 ppdiblc2 = -1.577008125e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.570251856e-05 lalpha0 = 2.076861164e-11 walpha0 = -1.041085477e-10 palpha0 = 9.834989220e-17   alpha1 = 0.0   beta0 = 1.884628103e+01 lbeta0 = 1.916771949e-06 wbeta0 = -2.046557818e-06 pbeta0 = 1.811031947e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.748119240e-01 lkt1 = 1.418405592e-08 wkt1 = 1.038536417e-08 pkt1 = -2.492946872e-14   kt2 = -2.522380507e-02 lkt2 = 6.114778183e-09 wkt2 = 2.354288428e-08 pkt2 = -2.852795610e-14   at = 8.908976513e+04 lat = -1.302394589e-02 wat = -2.153220828e-02 pat = 2.541490435e-8   ute = -2.892661567e-01 lute = -7.930879254e-07 wute = -1.266522246e-06 pute = 1.251797569e-12   ua1 = 7.784695216e-09 lua1 = -4.024033203e-15 wua1 = -8.718056636e-15 pua1 = 5.856326814e-21   ub1 = -1.020277097e-17 lub1 = 5.252768568e-24 wub1 = 1.328488438e-23 pub1 = -8.018143946e-30   uc1 = -2.677547992e-10 luc1 = 1.273787947e-16 wuc1 = 3.010743107e-16 puc1 = -1.552548433e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.45 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.975713447e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.222215947e-08 wvth0 = -8.432756760e-09 pvth0 = 2.539770520e-15   k1 = 2.201844036e-01 lk1 = 7.210549017e-08 wk1 = 2.460359286e-07 pk1 = -4.205919876e-14   k2 = 4.434774693e-02 lk2 = -2.218203883e-08 wk2 = -1.082118393e-07 pk2 = 1.955406125e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.567606882e+05 lvsat = 1.388583460e-03 wvsat = 2.255932024e-02 pvsat = -1.084068888e-8   ua = 7.434885225e-10 lua = -5.797126417e-16 wua = -3.800414833e-15 pua = 7.481244089e-22   ub = 3.959480243e-19 lub = 5.308454701e-25 wub = 3.743592548e-24 pub = -7.781420504e-31   uc = 2.500036568e-11 luc = 5.932603933e-18 wuc = 7.197581577e-17 puc = -1.868813680e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.263744916e-02 lu0 = -4.077411126e-09 wu0 = -2.790636689e-08 pu0 = 5.198452526e-15   a0 = 3.899166020e+00 la0 = -4.899508750e-07 wa0 = -5.510670775e-06 pa0 = 1.126288393e-12   keta = -1.565100049e-02 lketa = -5.050848466e-09 wketa = 6.164670755e-08 pketa = -7.931327272e-15   a1 = 0.0   a2 = 0.38689047   ags = 2.739243201e+00 lags = -5.524916573e-07 wags = -3.828325259e-06 pags = 7.721540631e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.668376836e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.619261185e-09 wvoff = -7.423891042e-08 pvoff = 1.429807848e-14   nfactor = {2.581872769e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.092218471e-08 wnfactor = -9.293858622e-08 pnfactor = -2.699028042e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.909525227e-06 lcit = -2.217607997e-12 wcit = -1.469440538e-11 pcit = 6.637389440e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.778153207e-02 leta0 = 6.551952601e-09 weta0 = 3.345811159e-08 peta0 = -1.067001265e-14   etab = 2.471163863e-02 letab = -1.119294093e-08 wetab = -2.956408414e-08 petab = 1.331181396e-14   dsub = 1.677296094e+00 ldsub = -3.059312593e-07 wdsub = -2.503538157e-07 pdsub = 1.130835668e-13   voffl = 0.0   minv = 0.0   pclm = 3.645531990e-01 lpclm = -4.867788084e-08 wpclm = -3.753249578e-07 ppclm = 2.200462658e-13   pdiblc1 = 0.39   pdiblc2 = 9.085031494e-03 lpdiblc2 = 2.789841470e-09 wpdiblc2 = -9.445252080e-09 ppdiblc2 = -1.608372209e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.075242670e-03 lalpha0 = 9.697550488e-10 walpha0 = 1.951235263e-09 palpha0 = -8.300386302e-16   alpha1 = 0.0   beta0 = 1.660735752e+01 lbeta0 = 2.928082504e-06 wbeta0 = 5.127530806e-06 pbeta0 = -1.429468014e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.213590357e-01 lkt1 = -9.960346477e-09 wkt1 = -8.030725277e-08 pkt1 = 1.603593289e-14   kt2 = -1.193464470e-02 lkt2 = 1.121308898e-10 wkt2 = -5.420034701e-08 pkt2 = 6.588272758e-15   at = 6.018430671e+04 lat = 3.250515771e-05 wat = 7.230701764e-02 pat = -1.697180480e-8   ute = -1.670714854e+00 lute = -1.690944562e-07 wute = 7.451106808e-07 pute = 3.431530341e-13   ua1 = -9.366839259e-10 lua1 = -8.462985196e-17 wua1 = 4.367088317e-15 pua1 = -5.416773522e-23   ub1 = 1.621384590e-18 lub1 = -8.814337818e-26 wub1 = -5.360904547e-24 pub1 = 4.040656844e-31   uc1 = 8.676665876e-11 luc1 = -3.275677521e-17 wuc1 = -1.868897125e-16 puc1 = 6.515606619e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.46 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.837134830e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.942709805e-08 wvth0 = 2.301997696e-07 pvth0 = -4.559121688e-14   k1 = 4.486605814e-01 lk1 = 2.602298748e-08 wk1 = -1.517359575e-07 pk1 = 3.816940180e-14   k2 = -5.733300750e-02 lk2 = -1.673539061e-09 wk2 = 4.105931719e-08 pk2 = -1.055318466e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.751939241e+05 lvsat = -2.329308053e-03 wvsat = -5.132270889e-02 pvsat = 4.060946991e-9   ua = -2.001180666e-09 lua = -2.612658968e-17 wua = -1.144326488e-16 pua = 4.680232146e-24   ub = 3.382016367e-18 lub = -7.142958431e-26 wub = 6.965009057e-25 pub = -1.635589016e-31   uc = 6.479536675e-11 luc = -2.093848808e-18 wuc = -3.820873140e-18 puc = -3.400323633e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.082161999e-02 lu0 = -1.694217462e-09 wu0 = 7.218461076e-09 pu0 = -1.886049651e-15   a0 = 4.235591648e+00 la0 = -5.578062421e-07 wa0 = 2.116235783e-07 pa0 = -2.786976715e-14   keta = 1.100620797e-01 lketa = -3.040654818e-08 wketa = 8.894756313e-09 pketa = 2.708477532e-15   a1 = 0.0   a2 = 0.38689047   ags = -2.255186821e+00 lags = 4.548599058e-07 wags = 3.221039076e-07 pags = -6.496674765e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.317407500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.468506731e-09 wvoff = -4.002357857e-08 pvoff = 7.397017128e-15   nfactor = {2.337176605e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.843180809e-08 wnfactor = -2.625797441e-06 pnfactor = 4.838746863e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.253401867e-05 lcit = 2.309142588e-12 wcit = 5.248001923e-11 pcit = -6.911356133e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.217794645e-01 leta0 = 2.752781557e-08 weta0 = -1.621154977e-08 peta0 = -6.518903068e-16   etab = -7.267203128e-02 letab = 8.448858368e-09 wetab = 1.404338962e-07 petab = -2.097592868e-14   dsub = -1.606983316e-01 ldsub = 6.478302642e-08 wdsub = 8.703758872e-07 pdsub = -1.129620106e-13   voffl = 0.0   minv = 0.0   pclm = 3.122316507e-02 lpclm = 1.855312034e-08 wpclm = 1.841465925e-06 ppclm = -2.270693712e-13   pdiblc1 = -7.452347020e-01 lpdiblc1 = 2.289711632e-07 wpdiblc1 = -2.036244958e-08 ppdiblc1 = 4.107004268e-15   pdiblc2 = 4.764832740e-02 lpdiblc2 = -4.988182498e-09 wpdiblc2 = -6.450838109e-08 ppdiblc2 = 9.497585597e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 6.682935824e-03 lalpha0 = -7.967257626e-10 walpha0 = -5.737767862e-09 palpha0 = 7.207948549e-16   alpha1 = 0.0   beta0 = 3.508042219e+01 lbeta0 = -7.978422756e-07 wbeta0 = -3.546216003e-06 pbeta0 = 3.199833485e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.149664578e-01 lkt1 = -1.124969746e-08 wkt1 = 9.409978771e-09 pkt1 = -2.059584127e-15   kt2 = 1.053874462e-02 lkt2 = -4.420639368e-09 wkt2 = -6.876173060e-08 pkt2 = 9.525231022e-15   at = 4.957125439e+04 lat = 2.173104745e-03 wat = -5.872897497e-02 pat = 9.457499732e-9   ute = -4.068638546e+00 lute = 3.145547629e-07 wute = 7.294463415e-06 pute = -9.778186656e-13   ua1 = -4.350235756e-09 lua1 = 6.038664843e-16 wua1 = 1.327342251e-14 pua1 = -1.850530809e-21   ub1 = 3.464068104e-18 lub1 = -4.598034296e-25 wub1 = -1.112816737e-23 pub1 = 1.567293759e-30   uc1 = -1.685469366e-10 luc1 = 1.873870040e-17 wuc1 = 2.781047102e-16 puc1 = -2.863098391e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.47 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.869708209e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.985607316e-08 wvth0 = -4.809899126e-07 pvth0 = 4.806890831e-14   k1 = 6.395864299e-01 lk1 = 8.790078641e-10 wk1 = 6.062178295e-07 pk1 = -6.164932217e-14   k2 = -1.338895597e-01 lk2 = 8.408576084e-09 wk2 = -1.469192108e-07 pk2 = 1.420264758e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.970696543e+05 lvsat = -5.210232347e-03 wvsat = -1.116784979e-01 pvsat = 1.200950262e-8   ua = -1.843181057e-09 lua = -4.693434823e-17 wua = 7.562800310e-17 pua = -2.034980540e-23   ub = 3.968631899e-18 lub = -1.486839168e-25 wub = -2.519898663e-24 pub = 2.600248396e-31   uc = 1.204025474e-10 luc = -9.417036468e-18 wuc = -1.301171174e-16 puc = 1.323226025e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.408265694e-02 lu0 = -2.123679723e-09 wu0 = -2.530271607e-08 pu0 = 2.396826773e-15   a0 = 0.0   keta = 6.592945011e-02 lketa = -2.459450152e-08 wketa = 1.293290822e-07 pketa = -1.315212101e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.033624482e+00 lags = 2.173990134e-08 wags = -7.515757844e-07 pags = 7.643149940e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.501734042e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.895995120e-09 wvoff = 7.087039828e-08 pvoff = -7.207165153e-15   nfactor = {1.301326928e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.548480312e-07 wnfactor = -6.271386468e-07 pnfactor = 2.206613164e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.194916667e-05 lcit = 2.232120504e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.147334562e-01 leta0 = -3.619753507e-09 weta0 = -9.289567844e-08 peta0 = 9.447026019e-15   etab = -3.738949304e-02 letab = 3.802324494e-09 wetab = -8.271622408e-08 petab = 8.411826408e-15   dsub = 5.726386546e-01 ldsub = -3.179378798e-08 wdsub = 5.540472764e-08 pdsub = -5.634383777e-15   voffl = 0.0   minv = 0.0   pclm = 1.859759373e-01 lpclm = -1.827045989e-09 wpclm = 5.147494575e-07 ppclm = -5.234744608e-14   pdiblc1 = 9.710826381e-01 lpdiblc1 = 2.940751122e-09 wpdiblc1 = 4.751238235e-08 ppdiblc1 = -4.831771724e-15   pdiblc2 = 2.312019524e-02 lpdiblc2 = -1.757950134e-09 wpdiblc2 = 3.340514497e-08 ppdiblc2 = -3.397136218e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.646109571e-03 lalpha0 = -1.334009293e-10 walpha0 = -1.161349454e-09 palpha0 = 1.181034327e-16   alpha1 = 0.0   beta0 = 3.261137501e+01 lbeta0 = -4.726811067e-07 wbeta0 = -4.901185600e-06 pbeta0 = 4.984260696e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.126897308e-01 lkt1 = -2.471903103e-08 wkt1 = -2.734456577e-08 pkt1 = 2.780805616e-15   kt2 = -6.159975487e-02 lkt2 = 5.079640322e-09 wkt2 = 1.565516368e-08 pkt2 = -1.592051870e-15   at = -5.164045768e+03 lat = 9.381470099e-03 wat = 5.743957910e-02 pat = -5.841317996e-9   ute = -1.736837580e+00 lute = 7.468234735e-09 wute = -5.724768741e-07 pute = 5.821803571e-14   ua1 = 5.134622809e-10 lua1 = -3.665822861e-17 wua1 = -3.416247751e-15 pua1 = 3.474153150e-22   ub1 = 1.493415477e-19 lub1 = -2.327051577e-26 wub1 = 3.392325253e-24 pub1 = -3.449825166e-31   uc1 = 1.763897157e-11 luc1 = -5.781052774e-18 wuc1 = 2.664671966e-16 puc1 = -2.709838156e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.48 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.49 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.50 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.164133052e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.875606883e-8   k1 = 6.067705922e-01 lk1 = -2.904914395e-7   k2 = -8.634485690e-02 lk2 = 1.150782937e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.545894796e+05 lvsat = -6.087170412e-1   ua = -8.523097748e-10 lua = -5.068737427e-16   ub = 2.210414102e-18 lub = 7.207334402e-25   uc = -6.060640140e-12 luc = 1.122725042e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.290174948e-02 lu0 = 8.748678201e-10   a0 = 1.977943329e+00 la0 = -2.180147316e-7   keta = 1.768528424e-01 lketa = -6.988684931e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.426975904e-01 lags = 3.760950596e-06 pags = -8.077935669e-28   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.035927842e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.624441498e-8   nfactor = {1.793948888e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.800957893e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378214013e-01 letab = 2.680094922e-7   dsub = 7.139466960e-01 ldsub = -6.083503888e-7   voffl = 0.0   minv = 0.0   pclm = 1.663039858e-01 lpclm = 1.331563707e-7   pdiblc1 = 0.39   pdiblc2 = 3.491130882e-03 lpdiblc2 = 1.611489017e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.896759563e-05 lalpha0 = 3.189117947e-10 palpha0 = -4.930380658e-32   alpha1 = 0.0   beta0 = 1.447755810e+01 lbeta0 = 1.310304963e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470030207e-01 lkt1 = -4.199458087e-8   kt2 = -3.565651056e-02 lkt2 = -2.795782473e-9   at = 6.706922666e+04 lat = -3.492992778e-2   ute = -1.240424282e+00 lute = 2.356169780e-7   ua1 = 1.882897412e-09 lua1 = 3.189120145e-16   ub1 = -1.048044516e-18 lub1 = -1.651632597e-24   uc1 = 1.342724329e-10 luc1 = -2.799951081e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.51 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.272507703e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.604642303e-9   k1 = 4.583582628e-01 lk1 = -8.358382679e-10   k2 = -2.242041396e-02 lk2 = -9.682721979e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.299730390e+03 lvsat = 7.689340581e-2   ua = -7.320202287e-10 lua = -7.416422484e-16   ub = 2.404845078e-18 lub = 3.412634777e-25   uc = 5.806214974e-11 luc = -1.287562416e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.793024204e-02 lu0 = -8.939215978e-9   a0 = 2.228395064e+00 la0 = -7.068201303e-7   keta = -2.466304804e-01 lketa = 1.276417906e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.249793801e+00 lags = 4.577236097e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.188380738e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.509740609e-9   nfactor = {8.611430018e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.404567944e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.475847500e-05 lcit = -9.287091865e-12 wcit = 6.462348536e-27   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.633067514e-04 leta0 = -1.235554702e-10   etab = -5.267331126e-04 letab = 5.217488210e-11   dsub = 2.399899413e-01 ldsub = 3.166686395e-7   voffl = 0.0   minv = 0.0   pclm = 2.560478239e-01 lpclm = -4.199622941e-8   pdiblc1 = 0.39   pdiblc2 = 8.945258225e-03 lpdiblc2 = 5.470097109e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.980734741e-04 lalpha0 = -1.437200758e-10   alpha1 = 0.0   beta0 = 2.158932331e+01 lbeta0 = -7.769469609e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675587881e-01 lkt1 = -1.875992557e-9   kt2 = -5.076961562e-02 lkt2 = 2.670038911e-8   at = 2.121024921e+04 lat = 5.457280922e-2   ute = -1.145205426e+00 lute = 4.977881240e-8   ua1 = 2.094550937e-09 lua1 = -9.417111151e-17   ub1 = -2.054850946e-18 lub1 = 3.133464795e-25   uc1 = 2.960755490e-11 luc1 = -7.572118907e-17 wuc1 = 6.162975822e-33   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.52 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.449224886e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.213443611e-9   k1 = 4.435587601e-01 lk1 = 1.324877441e-8   k2 = -2.204382508e-02 lk2 = -1.004111974e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.646641782e+04 lvsat = 6.436273521e-2   ua = -1.209922201e-09 lua = -2.868253308e-16   ub = 2.729363163e-18 lub = 3.242123834e-26 wub = -1.469367939e-39   uc = 3.348727667e-11 luc = 1.051215967e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.297005405e-02 lu0 = -4.218629868e-9   a0 = 1.944240793e+00 la0 = -4.363919315e-7   keta = -2.141504089e-01 lketa = 9.673066895e-8   a1 = 0.0   a2 = 0.38689047   ags = 3.089683441e+00 lags = -1.293290162e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.082137086e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.601414637e-9   nfactor = {1.133365243e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.813842489e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.623249313e-03 leta0 = 1.957379003e-09 peta0 = 3.944304526e-31   etab = -7.853050249e-04 letab = 2.982564782e-10   dsub = 1.867417334e-01 ldsub = 3.673446927e-7   voffl = 0.0   minv = 0.0   pclm = 1.099001673e-01 lpclm = 9.709176468e-8   pdiblc1 = 0.39   pdiblc2 = 2.133056769e-02 lpdiblc2 = -6.316939979e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.766084915e-05 lalpha0 = 8.062710091e-11 palpha0 = -1.232595164e-32   alpha1 = 0.0   beta0 = 1.760068882e+01 lbeta0 = 3.019016537e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.684911015e-01 lkt1 = -9.887145080e-10   kt2 = -1.089494863e-02 lkt2 = -1.124813209e-8   at = 7.598466223e+04 lat = 2.444274214e-3   ute = -1.060106943e+00 lute = -3.120898838e-8   ua1 = 2.478642633e-09 lua1 = -4.597092586e-16   ub1 = -2.117219565e-18 lub1 = 3.727023819e-25   uc1 = -8.451257089e-11 luc1 = 3.288636404e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.53 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.924389336e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.067638425e-8   k1 = 3.699287364e-01 lk1 = 4.650708796e-8   k2 = -2.151299859e-02 lk2 = -1.028089141e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.704909201e+05 lvsat = -5.209362345e-3   ua = -1.569550012e-09 lua = -1.243832468e-16   ub = 2.674402930e-18 lub = 5.724650092e-26   uc = 6.880685595e-11 luc = -5.441517696e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.565285543e-02 lu0 = -9.134878341e-10 wu0 = -1.323488980e-23   a0 = 5.452179876e-01 la0 = 1.955396745e-7   keta = 2.186890623e-02 lketa = -9.878075601e-9   a1 = 0.0   a2 = 0.38689047   ags = 4.092176022e-01 lags = -8.253714428e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.318676412e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.082948430e-9   nfactor = {2.525307752e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.734922266e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.661000000e-07 lcit = 1.822092461e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.582008429e-03 leta0 = 5.788510789e-11   etab = 6.718111913e-03 letab = -3.090999436e-09 wetab = 7.237830360e-25 petab = 7.395570986e-32   dsub = 1.524923775e+00 ldsub = -2.371054445e-7   voffl = 0.0   minv = 0.0   pclm = 1.361199546e-01 lpclm = 8.524841786e-8   pdiblc1 = 0.39   pdiblc2 = 3.336387468e-03 lpdiblc2 = 1.810941255e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.876664321e-04 lalpha0 = 4.645703727e-10 palpha0 = 2.465190329e-32   alpha1 = 0.0   beta0 = 1.972811587e+01 lbeta0 = 2.058068375e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702362710e-01 lkt1 = -2.004301707e-10   kt2 = -4.492248858e-02 lkt2 = 4.121937564e-9   at = 1.041923757e+05 lat = -1.029700891e-2   ute = -1.217219698e+00 lute = 3.975805749e-8   ua1 = 1.721247906e-09 lua1 = -1.175978474e-16 wua1 = -7.888609052e-31   ub1 = -1.641411537e-18 lub1 = 1.577822745e-25 wub1 = 7.346839693e-40   uc1 = -2.697963625e-11 luc1 = 6.899025125e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.54 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.238194875e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.717518506e-8   k1 = 3.563098429e-01 lk1 = 4.925395069e-8   k2 = -3.234316112e-02 lk2 = -8.096501780e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.439574911e+05 lvsat = 1.422976233e-4   ua = -2.070827570e-09 lua = -2.327806977e-17   ub = 3.805926257e-18 lub = -1.709760966e-25   uc = 6.246987672e-11 luc = -4.163380672e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.521497686e-02 lu0 = -2.842119918e-9   a0 = 4.364391664e+00 la0 = -5.747685602e-7   keta = 1.154756767e-01 lketa = -2.875809316e-08 pketa = -3.155443621e-30   a1 = 0.0   a2 = 0.38689047   ags = -2.059145393e+00 lags = 4.153193300e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.561002170e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.970537800e-9   nfactor = {7.390429982e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.129314468e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.940678571e-05 lcit = -1.897301645e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.316462661e-01 leta0 = 2.713105694e-08 weta0 = -2.646977960e-23 peta0 = 3.549874073e-30   etab = 1.279995733e-02 letab = -4.317677248e-9   dsub = 3.690367249e-01 ldsub = -3.968805937e-9   voffl = 0.0   minv = 0.0   pclm = 1.151990721e+00 lpclm = -1.196476363e-7   pdiblc1 = -7.576278571e-01 lpdiblc1 = 2.314708006e-7   pdiblc2 = 8.386726286e-03 lpdiblc2 = 7.923131668e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.190770166e-03 lalpha0 = -3.580298970e-10   alpha1 = 0.0   beta0 = 3.292209616e+01 lbeta0 = -6.030914792e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.092392821e-01 lkt1 = -1.250321784e-8   kt2 = -3.131156371e-02 lkt2 = 1.376682073e-9   at = 1.382716114e+04 lat = 7.929203033e-3   ute = 3.709754714e-01 lute = -2.805729672e-7   ua1 = 3.728339633e-09 lua1 = -5.224182132e-16   ub1 = -3.308845136e-18 lub1 = 4.940952943e-25   uc1 = 7.153517429e-13 luc1 = 1.313084522e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.55 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.168409367e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.674764481e-08 wvth0 = -2.014597077e-07 pvth0 = 2.653123621e-14   k1 = 1.082967320e+00 lk1 = -4.644320579e-08 wk1 = -1.222747085e-07 pk1 = 1.610296774e-14   k2 = -2.443757099e-01 lk2 = 1.982712473e-08 wk2 = 3.461395335e-08 pk2 = -4.558484587e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.564796732e+04 lvsat = 1.045527035e-02 wvsat = 1.042525908e-01 pvsat = -1.372954494e-8   ua = -3.538633562e-10 lua = -2.493936719e-16 wua = -2.371380552e-15 pua = 3.122989617e-22   ub = 1.806241172e-18 lub = 9.237243073e-26 wub = 1.032995798e-24 pub = -1.360403816e-31   uc = -5.272743913e-11 luc = 1.100752984e-17 wuc = 1.543423758e-16 puc = -2.032611918e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.507164607e-02 lu0 = -2.823243969e-09 wu0 = -2.692766477e-08 pu0 = 3.546238811e-15   a0 = 0.0   keta = 1.055683408e+00 lketa = -1.525787503e-07 wketa = -1.496876261e-06 pketa = 1.971311192e-13   a1 = 0.0   a2 = 0.38689047   ags = 5.679083539e-01 lags = 6.934948684e-08 wags = 1.361444215e-08 pags = -1.792953959e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.652825470e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.334930475e-08 wvoff = 2.599993243e-07 pvoff = -3.424061101e-14   nfactor = {-1.775089995e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.440301913e-07 wnfactor = 4.427537415e-06 pnfactor = -5.830845399e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.194916667e-05 lcit = 2.232120504e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.029811619e-01 leta0 = 2.335600604e-08 weta0 = 2.648181476e-07 peta0 = -3.487522595e-14   etab = -1.482476125e-01 letab = 1.689148246e-08 wetab = 9.942810045e-08 petab = -1.309418369e-14   dsub = 6.063595181e-01 ldsub = -3.522303120e-8   voffl = 0.0   minv = 0.0   pclm = 1.340050022e+00 lpclm = -1.444141060e-07 wpclm = -1.381440427e-06 ppclm = 1.819287970e-13   pdiblc1 = 7.409572600e-01 lpdiblc1 = 3.411463364e-08 wpdiblc1 = 4.256175835e-07 ppdiblc1 = -5.605170766e-14   pdiblc2 = 5.228140549e-02 lpdiblc2 = -4.988396611e-09 wpdiblc2 = -1.450788991e-08 ppdiblc2 = 1.910616562e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.699743888e-04 lalpha0 = 3.979380289e-11 walpha0 = 1.263999696e-09 palpha0 = -1.664624400e-16   alpha1 = 0.0   beta0 = 2.404909783e+01 lbeta0 = 5.654380360e-07 wbeta0 = 9.166978296e-06 pbeta0 = -1.207245207e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 1.952249366e-01 lkt1 = -6.576913313e-08 wkt1 = -5.332606809e-07 pkt1 = 7.022776537e-14   kt2 = -3.277992230e-02 lkt2 = 1.570057557e-09 wkt2 = -3.169697403e-08 pkt2 = 4.174332995e-15   at = -3.906762948e+04 lat = 1.489518248e-02 wat = 1.131445233e-01 pat = -1.490056799e-8   ute = -2.038135622e+00 lute = 3.669491824e-08 wute = -7.743213972e-08 pute = 1.019742564e-14   ua1 = -2.932869229e-09 lua1 = 3.548296879e-16 wua1 = 2.246212774e-15 pua1 = -2.958149913e-22   ub1 = 4.566825940e-18 lub1 = -5.430912081e-25 wub1 = -3.865778303e-24 pub1 = 5.091036736e-31   uc1 = 3.149858312e-10 luc1 = -4.007476626e-17 wuc1 = -2.220855876e-16 puc1 = 2.924756145e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.56 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.57 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.58 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.164133052e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.875606883e-8   k1 = 6.067705922e-01 lk1 = -2.904914395e-7   k2 = -8.634485690e-02 lk2 = 1.150782937e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.545894796e+05 lvsat = -6.087170412e-1   ua = -8.523097748e-10 lua = -5.068737427e-16   ub = 2.210414102e-18 lub = 7.207334402e-25   uc = -6.060640140e-12 luc = 1.122725042e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.290174948e-02 lu0 = 8.748678201e-10   a0 = 1.977943329e+00 la0 = -2.180147316e-7   keta = 1.768528424e-01 lketa = -6.988684931e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.426975904e-01 lags = 3.760950596e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.035927842e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.624441498e-8   nfactor = {1.793948888e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.800957893e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798762e-01 leta0 = -3.065720091e-7   etab = -1.378214012e-01 letab = 2.680094922e-7   dsub = 7.139466960e-01 ldsub = -6.083503888e-7   voffl = 0.0   minv = 0.0   pclm = 1.663039858e-01 lpclm = 1.331563707e-7   pdiblc1 = 0.39   pdiblc2 = 3.491130882e-03 lpdiblc2 = 1.611489017e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.896759563e-05 lalpha0 = 3.189117947e-10 palpha0 = -9.860761315e-32   alpha1 = 0.0   beta0 = 1.447755810e+01 lbeta0 = 1.310304963e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470030207e-01 lkt1 = -4.199458087e-8   kt2 = -3.565651056e-02 lkt2 = -2.795782473e-9   at = 6.706922665e+04 lat = -3.492992778e-2   ute = -1.240424282e+00 lute = 2.356169780e-7   ua1 = 1.882897412e-09 lua1 = 3.189120145e-16   ub1 = -1.048044516e-18 lub1 = -1.651632597e-24   uc1 = 1.342724329e-10 luc1 = -2.799951081e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.59 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.272507703e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.604642303e-9   k1 = 4.583582628e-01 lk1 = -8.358382679e-10   k2 = -2.242041396e-02 lk2 = -9.682721979e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.299730390e+03 lvsat = 7.689340581e-2   ua = -7.320202287e-10 lua = -7.416422484e-16   ub = 2.404845078e-18 lub = 3.412634777e-25   uc = 5.806214974e-11 luc = -1.287562416e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.793024204e-02 lu0 = -8.939215978e-9   a0 = 2.228395064e+00 la0 = -7.068201303e-7   keta = -2.466304804e-01 lketa = 1.276417906e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.249793801e+00 lags = 4.577236097e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.188380738e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.509740609e-9   nfactor = {8.611430018e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.404567944e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.475847500e-05 lcit = -9.287091865e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.633067514e-04 leta0 = -1.235554702e-10   etab = -5.267331126e-04 letab = 5.217488210e-11   dsub = 2.399899413e-01 ldsub = 3.166686395e-7   voffl = 0.0   minv = 0.0   pclm = 2.560478240e-01 lpclm = -4.199622941e-8   pdiblc1 = 0.39   pdiblc2 = 8.945258225e-03 lpdiblc2 = 5.470097109e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.980734741e-04 lalpha0 = -1.437200758e-10   alpha1 = 0.0   beta0 = 2.158932331e+01 lbeta0 = -7.769469609e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675587881e-01 lkt1 = -1.875992557e-9   kt2 = -5.076961562e-02 lkt2 = 2.670038911e-8   at = 2.121024921e+04 lat = 5.457280922e-2   ute = -1.145205426e+00 lute = 4.977881240e-8   ua1 = 2.094550937e-09 lua1 = -9.417111151e-17   ub1 = -2.054850947e-18 lub1 = 3.133464795e-25   uc1 = 2.960755490e-11 luc1 = -7.572118907e-17 wuc1 = 1.232595164e-32 puc1 = 2.350988702e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.60 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.449224886e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.213443611e-9   k1 = 4.435587601e-01 lk1 = 1.324877441e-8   k2 = -2.204382508e-02 lk2 = -1.004111974e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.646641782e+04 lvsat = 6.436273521e-2   ua = -1.209922201e-09 lua = -2.868253308e-16   ub = 2.729363163e-18 lub = 3.242123834e-26   uc = 3.348727667e-11 luc = 1.051215967e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.297005405e-02 lu0 = -4.218629868e-9   a0 = 1.944240793e+00 la0 = -4.363919315e-07 wa0 = -1.694065895e-21   keta = -2.141504089e-01 lketa = 9.673066895e-8   a1 = 0.0   a2 = 0.38689047   ags = 3.089683441e+00 lags = -1.293290162e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.082137086e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.601414637e-9   nfactor = {1.133365243e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.813842489e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.623249313e-03 leta0 = 1.957379003e-09 weta0 = -8.271806126e-25 peta0 = 7.888609052e-31   etab = -7.853050249e-04 letab = 2.982564782e-10   dsub = 1.867417334e-01 ldsub = 3.673446927e-7   voffl = 0.0   minv = 0.0   pclm = 1.099001673e-01 lpclm = 9.709176468e-8   pdiblc1 = 0.39   pdiblc2 = 2.133056769e-02 lpdiblc2 = -6.316939979e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.766084915e-05 lalpha0 = 8.062710091e-11   alpha1 = 0.0   beta0 = 1.760068882e+01 lbeta0 = 3.019016537e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.684911015e-01 lkt1 = -9.887145080e-10   kt2 = -1.089494863e-02 lkt2 = -1.124813209e-8   at = 7.598466223e+04 lat = 2.444274214e-3   ute = -1.060106943e+00 lute = -3.120898838e-8   ua1 = 2.478642633e-09 lua1 = -4.597092586e-16   ub1 = -2.117219565e-18 lub1 = 3.727023819e-25   uc1 = -8.451257089e-11 luc1 = 3.288636404e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.61 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.924389336e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.067638425e-8   k1 = 3.699287364e-01 lk1 = 4.650708796e-8   k2 = -2.151299859e-02 lk2 = -1.028089141e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.704909201e+05 lvsat = -5.209362345e-3   ua = -1.569550012e-09 lua = -1.243832468e-16   ub = 2.674402930e-18 lub = 5.724650092e-26   uc = 6.880685595e-11 luc = -5.441517696e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.565285543e-02 lu0 = -9.134878341e-10   a0 = 5.452179876e-01 la0 = 1.955396745e-7   keta = 2.186890623e-02 lketa = -9.878075601e-9   a1 = 0.0   a2 = 0.38689047   ags = 4.092176022e-01 lags = -8.253714428e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.318676412e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.082948430e-9   nfactor = {2.525307752e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.734922266e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.661000000e-07 lcit = 1.822092461e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.582008429e-03 leta0 = 5.788510789e-11   etab = 6.718111913e-03 letab = -3.090999436e-09 wetab = 2.895132144e-24 petab = 1.479114197e-31   dsub = 1.524923775e+00 ldsub = -2.371054445e-7   voffl = 0.0   minv = 0.0   pclm = 1.361199546e-01 lpclm = 8.524841786e-8   pdiblc1 = 0.39   pdiblc2 = 3.336387468e-03 lpdiblc2 = 1.810941255e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.876664321e-04 lalpha0 = 4.645703727e-10 walpha0 = -2.067951531e-25 palpha0 = -4.930380658e-32   alpha1 = 0.0   beta0 = 1.972811587e+01 lbeta0 = 2.058068375e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702362710e-01 lkt1 = -2.004301707e-10   kt2 = -4.492248858e-02 lkt2 = 4.121937564e-9   at = 1.041923757e+05 lat = -1.029700891e-2   ute = -1.217219698e+00 lute = 3.975805749e-8   ua1 = 1.721247906e-09 lua1 = -1.175978474e-16   ub1 = -1.641411537e-18 lub1 = 1.577822745e-25   uc1 = -2.697963625e-11 luc1 = 6.899025125e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.62 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.238194875e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.717518506e-8   k1 = 3.563098429e-01 lk1 = 4.925395069e-8   k2 = -3.234316112e-02 lk2 = -8.096501780e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.439574911e+05 lvsat = 1.422976233e-4   ua = -2.070827570e-09 lua = -2.327806977e-17   ub = 3.805926257e-18 lub = -1.709760966e-25   uc = 6.246987672e-11 luc = -4.163380672e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.521497686e-02 lu0 = -2.842119918e-9   a0 = 4.364391664e+00 la0 = -5.747685602e-7   keta = 1.154756767e-01 lketa = -2.875809316e-08 pketa = -1.262177448e-29   a1 = 0.0   a2 = 0.38689047   ags = -2.059145393e+00 lags = 4.153193300e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.561002170e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.970537800e-9   nfactor = {7.390429982e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.129314468e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.940678571e-05 lcit = -1.897301645e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.316462661e-01 leta0 = 2.713105694e-08 weta0 = -3.308722450e-23 peta0 = -8.677469957e-30   etab = 1.279995733e-02 letab = -4.317677248e-9   dsub = 3.690367249e-01 ldsub = -3.968805937e-9   voffl = 0.0   minv = 0.0   pclm = 1.151990721e+00 lpclm = -1.196476363e-7   pdiblc1 = -7.576278571e-01 lpdiblc1 = 2.314708006e-07 ppdiblc1 = -1.009741959e-28   pdiblc2 = 8.386726286e-03 lpdiblc2 = 7.923131668e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.190770166e-03 lalpha0 = -3.580298970e-10 palpha0 = 3.944304526e-31   alpha1 = 0.0   beta0 = 3.292209616e+01 lbeta0 = -6.030914792e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.092392821e-01 lkt1 = -1.250321784e-8   kt2 = -3.131156371e-02 lkt2 = 1.376682073e-9   at = 1.382716114e+04 lat = 7.929203033e-3   ute = 3.709754714e-01 lute = -2.805729672e-7   ua1 = 3.728339633e-09 lua1 = -5.224182132e-16   ub1 = -3.308845136e-18 lub1 = 4.940952943e-25 wub1 = -1.469367939e-39 pub1 = -3.503246161e-46   uc1 = 7.153517429e-13 luc1 = 1.313084522e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.63 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.900206672e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.752264400e-07 wvth0 = 2.000157250e-06 pvth0 = -2.634107090e-13   k1 = 1.939364397e+00 lk1 = -1.592264189e-07 wk1 = -9.727112620e-07 pk1 = 1.281012097e-13   k2 = -5.050046722e-01 lk2 = 5.415065592e-08 wk2 = 2.934289381e-07 pk2 = -3.864312400e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.754672951e+05 lvsat = -1.717688602e-02 wvsat = -1.041063945e-01 pvsat = 1.371029163e-8   ua = -6.408943064e-09 lua = 5.480300503e-16 wua = 3.641555802e-15 pua = -4.795746913e-22   ub = 5.130120411e-18 lub = -3.453658457e-25 wub = -2.267749242e-24 pub = 2.986512364e-31   uc = 1.798595757e-11 luc = 1.694929062e-18 wuc = 8.412114431e-17 puc = -1.107833410e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -4.216838379e-02 lu0 = 7.348881764e-09 wu0 = 4.977477449e-08 pu0 = -6.555088927e-15   a0 = 0.0   keta = -2.354440852e+00 lketa = 2.965175641e-07 wketa = 1.889513534e-06 pketa = -2.488394849e-13   a1 = 0.0   a2 = 0.38689047   ags = 5.339654651e-01 lags = 7.381959557e-08 wags = 4.732108842e-08 pags = -6.231950740e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {5.316218490e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.159901967e-08 wvoff = -5.313586171e-07 pvoff = 6.997727307e-14   nfactor = {1.288244746e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.286294204e-06 wnfactor = -1.012798358e-05 pnfactor = 1.333804798e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.194916667e-05 lcit = 2.232120504e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.688740326e-01 leta0 = 3.203376765e-08 weta0 = 3.302524039e-07 peta0 = -4.349259033e-14   etab = 1.215020041e-01 letab = -1.863319329e-08 wetab = -1.684440587e-07 petab = 2.218324031e-14   dsub = 6.070439528e-01 ldsub = -3.531316783e-08 wdsub = -6.796710404e-10 pdsub = 8.950927767e-17   voffl = 0.0   minv = 0.0   pclm = -5.742631854e-02 lpclm = 3.962654067e-08 wpclm = 6.309478457e-09 ppclm = -8.309267653e-16   pdiblc1 = 2.052361131e+00 lpdiblc1 = -1.385906992e-07 wpdiblc1 = -8.766589168e-07 ppdiblc1 = 1.154515960e-13   pdiblc2 = 2.355772401e-01 lpdiblc2 = -2.912754155e-08 wpdiblc2 = -1.965279855e-07 ppdiblc2 = 2.588175305e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.701707651e-03 lalpha0 = 2.862849692e-10 walpha0 = 3.122654829e-09 palpha0 = -4.112380277e-16   alpha1 = 0.0   beta0 = -7.766276344e+01 lbeta0 = 1.396038161e-05 wbeta0 = 1.101709250e-04 pbeta0 = -1.450895997e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -7.688830991e-01 lkt1 = 6.119907464e-08 wkt1 = 4.241371629e-07 pkt1 = -5.585674367e-14   kt2 = -2.688310868e-01 lkt2 = 3.265681567e-08 wkt2 = 2.027112744e-07 pkt2 = -2.669606128e-14   at = 1.396776411e+05 lat = -8.644675930e-03 wat = -6.435668026e-02 pat = 8.475453006e-9   ute = -3.346257424e+00 lute = 2.089680190e-07 wute = 1.221585135e-06 pute = -1.608766543e-13   ua1 = -2.723158409e-09 lua1 = 3.272118214e-16 wua1 = 2.037961541e-15 pua1 = -2.683893452e-22   ub1 = 2.044853945e-19 lub1 = 3.140723012e-26 wub1 = 4.662003526e-25 pub1 = -6.139625544e-32   uc1 = 6.582878939e-10 luc1 = -8.528593142e-17 wuc1 = -5.629982679e-16 puc1 = 7.414405690e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.64 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.65 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.66 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.164133052e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.875606883e-8   k1 = 6.067705922e-01 lk1 = -2.904914395e-7   k2 = -8.634485690e-02 lk2 = 1.150782937e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.545894796e+05 lvsat = -6.087170412e-1   ua = -8.523097748e-10 lua = -5.068737427e-16   ub = 2.210414102e-18 lub = 7.207334402e-25   uc = -6.060640140e-12 luc = 1.122725042e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.290174948e-02 lu0 = 8.748678201e-10   a0 = 1.977943329e+00 la0 = -2.180147316e-7   keta = 1.768528424e-01 lketa = -6.988684931e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.426975904e-01 lags = 3.760950596e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.035927842e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.624441498e-8   nfactor = {1.793948888e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.800957893e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378214013e-01 letab = 2.680094922e-7   dsub = 7.139466960e-01 ldsub = -6.083503888e-7   voffl = 0.0   minv = 0.0   pclm = 1.663039858e-01 lpclm = 1.331563707e-7   pdiblc1 = 0.39   pdiblc2 = 3.491130882e-03 lpdiblc2 = 1.611489017e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.896759563e-05 lalpha0 = 3.189117947e-10 palpha0 = -4.930380658e-32   alpha1 = 0.0   beta0 = 1.447755810e+01 lbeta0 = 1.310304963e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470030207e-01 lkt1 = -4.199458087e-8   kt2 = -3.565651056e-02 lkt2 = -2.795782473e-9   at = 6.706922666e+04 lat = -3.492992778e-2   ute = -1.240424282e+00 lute = 2.356169780e-7   ua1 = 1.882897412e-09 lua1 = 3.189120145e-16   ub1 = -1.048044516e-18 lub1 = -1.651632597e-24   uc1 = 1.342724329e-10 luc1 = -2.799951081e-16 wuc1 = 4.930380658e-32   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.67 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.272507703e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.604642303e-9   k1 = 4.583582628e-01 lk1 = -8.358382679e-10   k2 = -2.242041396e-02 lk2 = -9.682721979e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.299730390e+03 lvsat = 7.689340581e-2   ua = -7.320202287e-10 lua = -7.416422484e-16   ub = 2.404845078e-18 lub = 3.412634777e-25   uc = 5.806214974e-11 luc = -1.287562416e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.793024204e-02 lu0 = -8.939215978e-9   a0 = 2.228395064e+00 la0 = -7.068201303e-7   keta = -2.466304804e-01 lketa = 1.276417906e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.249793801e+00 lags = 4.577236097e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.188380738e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.509740609e-9   nfactor = {8.611430018e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.404567944e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.475847500e-05 lcit = -9.287091865e-12 wcit = -6.462348536e-27   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.633067514e-04 leta0 = -1.235554702e-10   etab = -5.267331125e-04 letab = 5.217488210e-11   dsub = 2.399899413e-01 ldsub = 3.166686395e-7   voffl = 0.0   minv = 0.0   pclm = 2.560478239e-01 lpclm = -4.199622941e-8   pdiblc1 = 0.39   pdiblc2 = 8.945258225e-03 lpdiblc2 = 5.470097109e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.980734741e-04 lalpha0 = -1.437200758e-10   alpha1 = 0.0   beta0 = 2.158932331e+01 lbeta0 = -7.769469609e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675587881e-01 lkt1 = -1.875992557e-9   kt2 = -5.076961563e-02 lkt2 = 2.670038911e-8   at = 2.121024920e+04 lat = 5.457280922e-2   ute = -1.145205426e+00 lute = 4.977881240e-8   ua1 = 2.094550936e-09 lua1 = -9.417111151e-17   ub1 = -2.054850946e-18 lub1 = 3.133464795e-25   uc1 = 2.960755490e-11 luc1 = -7.572118907e-17 wuc1 = -6.162975822e-33 puc1 = 1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.68 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.449224886e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.213443611e-9   k1 = 4.435587601e-01 lk1 = 1.324877441e-8   k2 = -2.204382508e-02 lk2 = -1.004111974e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.646641782e+04 lvsat = 6.436273521e-2   ua = -1.209922201e-09 lua = -2.868253308e-16   ub = 2.729363163e-18 lub = 3.242123834e-26   uc = 3.348727667e-11 luc = 1.051215967e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.297005405e-02 lu0 = -4.218629868e-9   a0 = 1.944240793e+00 la0 = -4.363919315e-7   keta = -2.141504089e-01 lketa = 9.673066895e-8   a1 = 0.0   a2 = 0.38689047   ags = 3.089683441e+00 lags = -1.293290162e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.082137086e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.601414637e-9   nfactor = {1.133365243e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.813842489e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.623249313e-03 leta0 = 1.957379003e-09 peta0 = 1.972152263e-31   etab = -7.853050249e-04 letab = 2.982564782e-10   dsub = 1.867417334e-01 ldsub = 3.673446927e-7   voffl = 0.0   minv = 0.0   pclm = 1.099001673e-01 lpclm = 9.709176468e-8   pdiblc1 = 0.39   pdiblc2 = 2.133056769e-02 lpdiblc2 = -6.316939979e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.766084915e-05 lalpha0 = 8.062710091e-11 palpha0 = 1.232595164e-32   alpha1 = 0.0   beta0 = 1.760068882e+01 lbeta0 = 3.019016537e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.684911015e-01 lkt1 = -9.887145080e-10   kt2 = -1.089494863e-02 lkt2 = -1.124813209e-8   at = 7.598466223e+04 lat = 2.444274214e-3   ute = -1.060106943e+00 lute = -3.120898838e-8   ua1 = 2.478642633e-09 lua1 = -4.597092586e-16   ub1 = -2.117219565e-18 lub1 = 3.727023819e-25   uc1 = -8.451257089e-11 luc1 = 3.288636404e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.69 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.924389336e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.067638425e-8   k1 = 3.699287364e-01 lk1 = 4.650708796e-8   k2 = -2.151299859e-02 lk2 = -1.028089141e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.704909201e+05 lvsat = -5.209362345e-3   ua = -1.569550012e-09 lua = -1.243832468e-16   ub = 2.674402930e-18 lub = 5.724650092e-26   uc = 6.880685595e-11 luc = -5.441517696e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.565285543e-02 lu0 = -9.134878341e-10 wu0 = 1.323488980e-23   a0 = 5.452179876e-01 la0 = 1.955396745e-7   keta = 2.186890623e-02 lketa = -9.878075601e-9   a1 = 0.0   a2 = 0.38689047   ags = 4.092176022e-01 lags = -8.253714428e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.318676412e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.082948430e-9   nfactor = {2.525307752e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.734922266e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.661000000e-07 lcit = 1.822092460e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.582008429e-03 leta0 = 5.788510789e-11   etab = 6.718111913e-03 letab = -3.090999436e-09 wetab = 1.447566072e-24 petab = -7.642090019e-31   dsub = 1.524923775e+00 ldsub = -2.371054445e-7   voffl = 0.0   minv = 0.0   pclm = 1.361199546e-01 lpclm = 8.524841786e-8   pdiblc1 = 0.39   pdiblc2 = 3.336387468e-03 lpdiblc2 = 1.810941255e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.876664321e-04 lalpha0 = 4.645703727e-10 walpha0 = 1.033975766e-25 palpha0 = -4.930380658e-32   alpha1 = 0.0   beta0 = 1.972811587e+01 lbeta0 = 2.058068375e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702362710e-01 lkt1 = -2.004301707e-10   kt2 = -4.492248858e-02 lkt2 = 4.121937564e-9   at = 1.041923757e+05 lat = -1.029700891e-2   ute = -1.217219698e+00 lute = 3.975805749e-8   ua1 = 1.721247906e-09 lua1 = -1.175978474e-16 wua1 = 7.888609052e-31   ub1 = -1.641411537e-18 lub1 = 1.577822745e-25   uc1 = -2.697963625e-11 luc1 = 6.899025125e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.70 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.238194875e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.717518506e-8   k1 = 3.563098429e-01 lk1 = 4.925395069e-8   k2 = -3.234316112e-02 lk2 = -8.096501780e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.439574911e+05 lvsat = 1.422976233e-4   ua = -2.070827570e-09 lua = -2.327806977e-17   ub = 3.805926257e-18 lub = -1.709760966e-25   uc = 6.246987672e-11 luc = -4.163380672e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.521497686e-02 lu0 = -2.842119918e-9   a0 = 4.364391664e+00 la0 = -5.747685602e-7   keta = 1.154756767e-01 lketa = -2.875809316e-08 wketa = -2.646977960e-23   a1 = 0.0   a2 = 0.38689047   ags = -2.059145393e+00 lags = 4.153193300e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.561002170e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.970537800e-9   nfactor = {7.390429982e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.129314468e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.940678571e-05 lcit = -1.897301645e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.316462661e-01 leta0 = 2.713105694e-08 weta0 = 2.316105715e-23 peta0 = 2.366582716e-30   etab = 1.279995733e-02 letab = -4.317677248e-9   dsub = 3.690367249e-01 ldsub = -3.968805937e-9   voffl = 0.0   minv = 0.0   pclm = 1.151990721e+00 lpclm = -1.196476363e-7   pdiblc1 = -7.576278571e-01 lpdiblc1 = 2.314708006e-7   pdiblc2 = 8.386726286e-03 lpdiblc2 = 7.923131668e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.190770166e-03 lalpha0 = -3.580298970e-10   alpha1 = 0.0   beta0 = 3.292209616e+01 lbeta0 = -6.030914792e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.092392821e-01 lkt1 = -1.250321784e-8   kt2 = -3.131156371e-02 lkt2 = 1.376682073e-9   at = 1.382716114e+04 lat = 7.929203033e-3   ute = 3.709754714e-01 lute = -2.805729672e-7   ua1 = 3.728339633e-09 lua1 = -5.224182132e-16 pua1 = -1.880790961e-37   ub1 = -3.308845136e-18 lub1 = 4.940952943e-25 pub1 = -1.751623080e-46   uc1 = 7.153517429e-13 luc1 = 1.313084522e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.71 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.532955044e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.471802911e-08 wvth0 = 3.959579659e-08 pvth0 = -5.214568433e-15   k1 = 7.716998650e-01 lk1 = -5.450838271e-9   k2 = -1.406952704e-01 lk2 = 6.172929254e-09 wk2 = -1.005536595e-08 pk2 = 1.324241419e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.032480418e+04 lvsat = 9.839354324e-03 wvsat = 6.678550613e-02 pvsat = -8.795317230e-9   ua = -2.041142479e-09 lua = -2.718744774e-17 wua = 3.003202631e-18 pua = -3.955067705e-25   ub = 3.132179474e-18 lub = -8.224701404e-26 wub = -6.033845239e-25 pub = 7.946272487e-32   uc = 1.189668760e-10 luc = -1.160375299e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.171108965e-02 lu0 = -1.063725490e-09 wu0 = -3.439382061e-09 pu0 = 4.529494205e-16   a0 = 0.0   keta = 3.940477007e-01 lketa = -6.544463587e-08 wketa = -4.000873696e-07 pketa = 5.268950613e-14   a1 = 0.0   a2 = 0.38689047   ags = 5.907707667e-01 lags = 6.633862138e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.062350121e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.403539648e-09 wvoff = 1.662487171e-12 pvoff = -2.189412480e-19   nfactor = {3.370868675e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.366683571e-08 wnfactor = -2.204457988e-06 pnfactor = 2.903160948e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.194916667e-05 lcit = 2.232120504e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.275683998e-01 leta0 = -2.017571849e-8   etab = -8.070204224e-02 letab = 7.996068586e-9   dsub = 6.062280604e-01 ldsub = -3.520571887e-8   voffl = 0.0   minv = 0.0   pclm = -2.256014960e-01 lpclm = 6.177437066e-08 wpclm = 1.464061283e-07 ppclm = -1.928095506e-14   pdiblc1 = 1.0   pdiblc2 = -7.882223995e-03 lpdiblc2 = 2.934852574e-09 wpdiblc2 = 6.283486457e-09 ppdiblc2 = -8.275037490e-16   pdiblcb = 0.0   drout = -2.275190404e+01 ldrout = 3.456533350e-06 wdrout = 2.186438773e-05 pdrout = -2.879430542e-12   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.019554343e-03 lalpha0 = -2.037866292e-10 walpha0 = 2.269473750e-11 palpha0 = -2.988783455e-18   alpha1 = 0.0   beta0 = 4.833360039e+01 lbeta0 = -2.632709528e-06 wbeta0 = 5.210914089e-06 pbeta0 = -6.862513310e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.099522915e-01 lkt1 = 1.392968193e-08 wkt1 = 1.251334430e-07 pkt1 = -1.647944877e-14   kt2 = -2.549190217e-02 lkt2 = 6.102617458e-10   at = 1.111129041e+05 lat = -4.882842888e-03 wat = -4.056111173e-02 pat = 5.341695609e-9   ute = -1.879839083e+00 lute = 1.584805558e-8   ua1 = -2.767434217e-10 lua1 = 5.031199616e-18   ub1 = 7.641228100e-19 lub1 = -4.229421931e-26   uc1 = -1.754792183e-11 luc1 = 3.718266336e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.72 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.73 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4236902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057223608   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.805772e-10   ub = 2.3928e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03312314   a0 = 1.9227734   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.5090334   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5459298+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.74 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.164133052e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.875606883e-8   k1 = 6.067705922e-01 lk1 = -2.904914395e-7   k2 = -8.634485690e-02 lk2 = 1.150782937e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.545894796e+05 lvsat = -6.087170412e-1   ua = -8.523097748e-10 lua = -5.068737427e-16   ub = 2.210414102e-18 lub = 7.207334402e-25   uc = -6.060640140e-12 luc = 1.122725042e-16 puc = 4.701977403e-38   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.290174948e-02 lu0 = 8.748678201e-10   a0 = 1.977943329e+00 la0 = -2.180147316e-7   keta = 1.768528424e-01 lketa = -6.988684931e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.426975904e-01 lags = 3.760950596e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.035927842e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.624441498e-8   nfactor = {1.793948888e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.800957893e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.575798763e-01 leta0 = -3.065720091e-7   etab = -1.378214013e-01 letab = 2.680094922e-7   dsub = 7.139466960e-01 ldsub = -6.083503888e-7   voffl = 0.0   minv = 0.0   pclm = 1.663039858e-01 lpclm = 1.331563707e-7   pdiblc1 = 0.39   pdiblc2 = 3.491130882e-03 lpdiblc2 = 1.611489017e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.896759563e-05 lalpha0 = 3.189117947e-10 palpha0 = -9.860761315e-32   alpha1 = 0.0   beta0 = 1.447755810e+01 lbeta0 = 1.310304963e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470030207e-01 lkt1 = -4.199458087e-8   kt2 = -3.565651056e-02 lkt2 = -2.795782473e-9   at = 6.706922666e+04 lat = -3.492992778e-2   ute = -1.240424282e+00 lute = 2.356169780e-7   ua1 = 1.882897412e-09 lua1 = 3.189120145e-16   ub1 = -1.048044516e-18 lub1 = -1.651632597e-24   uc1 = 1.342724329e-10 luc1 = -2.799951081e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.75 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.698113917e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.148782903e-07 wvth0 = 9.966542423e-08 pvth0 = -1.945165101e-13   k1 = 5.858951043e-01 lk1 = -2.497488542e-07 wk1 = -8.073592216e-08 pk1 = 1.575718956e-13   k2 = -7.128063356e-02 lk2 = 8.567752430e-08 wk2 = 3.093047341e-08 pk2 = -6.036685030e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.674035201e+04 lvsat = -7.889438198e-03 wvsat = -2.749965111e-02 pvsat = 5.367093157e-8   ua = 1.116102705e-09 lua = -4.348614537e-15 wua = -1.169935742e-15 pua = 2.283357738e-21   ub = 2.749613739e-18 lub = -3.316197945e-25 wub = -2.182523533e-25 pub = 4.259620266e-31   uc = -5.300572908e-11 luc = 2.038949996e-16 wuc = 7.031041001e-17 puc = -1.372244757e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.788355507e-02 lu0 = -8.691589724e-08 wu0 = -2.529204528e-08 pu0 = 4.936235830e-14   a0 = 2.653906432e+00 la0 = -1.537288541e-06 wa0 = -2.693657167e-07 pa0 = 5.257197224e-13   keta = -3.470635897e-01 lketa = 3.236565879e-07 wketa = 6.357817553e-08 pketa = -1.240852073e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.410291537e+00 lags = 1.444809805e-07 wags = -1.016014869e-07 pags = 1.982951140e-13   b0 = 5.536339262e-07 lb0 = -1.080524566e-12 wb0 = -3.504724207e-13 pb0 = 6.840152710e-19   b1 = 6.005888453e-09 lb1 = -1.172166246e-14 wb1 = -3.801967626e-15 pb1 = 7.420281207e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.050111746e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.716933506e-07 wvoff = 5.455101973e-08 pvoff = -1.064669525e-13   nfactor = {-3.721577973e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.784530407e-06 wnfactor = 2.901045686e-06 pnfactor = -5.661956360e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 4.347005571e-05 lcit = -6.532334038e-11 wcit = -1.817557905e-11 pcit = 3.547318676e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.557514354e-03 leta0 = 4.015640477e-09 weta0 = 1.342564593e-09 peta0 = -2.620276603e-15   etab = 2.183123298e-03 letab = -5.236638325e-09 wetab = -1.715447502e-09 petab = 3.348030313e-15   dsub = -1.555814175e+00 ldsub = 3.821530555e-06 wdsub = 1.136815838e-06 pdsub = -2.218717787e-12   voffl = 0.0   minv = 0.0   pclm = 4.418691743e-01 lpclm = -4.046628298e-07 wpclm = -1.176323476e-07 ppclm = 2.295824647e-13   pdiblc1 = 0.39   pdiblc2 = -9.476091959e-03 lpdiblc2 = 4.142295416e-08 wpdiblc2 = 1.166145152e-08 ppdiblc2 = -2.275959663e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.355168454e-04 lalpha0 = -6.071371165e-10 walpha0 = -1.503111518e-10 palpha0 = 2.933615234e-16   alpha1 = 0.0   beta0 = 2.806702917e+01 lbeta0 = -1.341945310e-05 wbeta0 = -4.100646917e-06 pbeta0 = 8.003212085e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.872237852e-01 lkt1 = -1.586654159e-07 wkt1 = -5.085527019e-08 pkt1 = 9.925397656e-14   kt2 = -1.026686689e-01 lkt2 = 1.279915119e-07 wkt2 = 3.285417670e-08 pkt2 = -6.412133239e-14   at = 5.847213865e+04 lat = -1.815103411e-02 wat = -2.358826650e-02 pat = 4.603710178e-8   ute = -9.356108868e-01 lute = -3.592858018e-07 wute = -1.326817271e-07 pute = 2.589542634e-13   ua1 = 2.739987271e-09 lua1 = -1.353865978e-15 wua1 = -4.085870171e-16 pua1 = 7.974372384e-22   ub1 = -3.036212775e-18 lub1 = 2.228665454e-24 wub1 = 6.212412920e-25 pub1 = -1.212473523e-30   uc1 = 5.337082621e-10 luc1 = -1.059572019e-15 wuc1 = -3.191159117e-16 puc1 = 6.228169292e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.76 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {7.598012458e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.514426038e-07 wvth0 = -1.993308485e-07 pvth0 = 9.003674759e-14   k1 = 1.884850771e-01 lk1 = 1.284642817e-07 wk1 = 1.614718443e-07 pk1 = -7.293602472e-14   k2 = 7.567661410e-02 lk2 = -5.418095352e-08 wk2 = -6.186094682e-08 pk2 = 2.794228037e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -7.041482541e+04 lvsat = 1.036065584e-01 wvsat = 5.499930222e-02 pvsat = -2.484290981e-8   ua = -4.906168068e-09 lua = 1.382750446e-15 wua = 2.339871484e-15 pua = -1.056908250e-21   ub = 2.039825841e-18 lub = 3.438817992e-25 wub = 4.365047065e-25 pub = -1.971669934e-31   uc = 2.556230343e-10 luc = -8.982545138e-17 wuc = -1.406208200e-16 puc = 6.351772130e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -4.693657199e-02 lu0 = 3.187479358e-08 wu0 = 5.058409055e-08 pu0 = -2.284858078e-14   a0 = 1.093218056e+00 la0 = -5.198921636e-08 wa0 = 5.387314334e-07 pa0 = -2.433422948e-13   keta = -1.328419025e-02 lketa = 6.000402313e-09 wketa = -1.271563511e-07 pketa = 5.743588799e-14   a1 = 0.0   a2 = 0.38689047   ags = 2.768687969e+00 lags = -1.148298112e-06 wags = 2.032029738e-07 pags = -9.178576726e-14   b0 = -1.107267852e-06 lb0 = 5.001473526e-13 wb0 = 7.009448413e-13 pb0 = -3.166132801e-19   b1 = -1.201177691e-08 lb1 = 5.425659570e-15 wb1 = 7.603935253e-15 pb1 = -3.434659534e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {6.413249298e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.444933217e-08 wvoff = -1.091020395e-07 pvoff = 4.928084572e-14   nfactor = {1.029880719e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.558600052e-06 wnfactor = -5.802091371e-06 pnfactor = 2.620775662e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -5.242316142e-05 lcit = 2.593775490e-11 wcit = 3.635115811e-11 pcit = -1.641963636e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.618392898e-03 leta0 = 4.145042493e-11 weta0 = -2.685129185e-09 peta0 = 1.212859427e-15   etab = -6.205017846e-03 letab = 2.746313661e-09 wetab = 3.430895004e-09 petab = -1.549718119e-15   dsub = 3.778349967e+00 ldsub = -1.254966788e-06 wdsub = -2.273631676e-06 pdsub = 1.026988060e-12   voffl = 0.0   minv = 0.0   pclm = -2.617425334e-01 lpclm = 2.649609144e-07 wpclm = 2.352646953e-07 ppclm = -1.062678865e-13   pdiblc1 = 0.39   pdiblc2 = 5.817326805e-02 lpdiblc2 = -2.295860352e-08 wpdiblc2 = -2.332290304e-08 ppdiblc2 = 1.053483869e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.125475919e-04 lalpha0 = 2.951310682e-10 walpha0 = 3.006223036e-10 palpha0 = -1.357895914e-16   alpha1 = 0.0   beta0 = 4.645277104e+00 lbeta0 = 8.870911233e-06 wbeta0 = 8.201293834e-06 pbeta0 = -3.704483418e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.291611072e-01 lkt1 = 7.158512370e-08 wkt1 = 1.017105404e-07 pkt1 = -4.594214254e-14   kt2 = 9.290315796e-02 lkt2 = -5.813321785e-08 wkt2 = -6.570835339e-08 pkt2 = 2.968013469e-14   at = 1.460883336e+03 lat = 3.610629252e-02 wat = 4.717653299e-02 pat = -2.130940407e-8   ute = -1.479296021e+00 lute = 1.581366224e-07 wute = 2.653634542e-07 pute = -1.198633454e-13   ua1 = 1.187769964e-09 lua1 = 1.233714715e-16 wua1 = 8.171740342e-16 pua1 = -3.691134254e-22   ub1 = -1.544959076e-19 lub1 = -5.138500805e-25 wub1 = -1.242482584e-24 pub1 = 5.612231708e-31   uc1 = -1.092713985e-09 luc1 = 4.882859019e-16 wuc1 = 6.382318233e-16 puc1 = -2.882861234e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.77 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.924389336e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.067638425e-8   k1 = 3.699287364e-01 lk1 = 4.650708796e-8   k2 = -2.151299859e-02 lk2 = -1.028089141e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.704909201e+05 lvsat = -5.209362345e-3   ua = -1.569550012e-09 lua = -1.243832468e-16   ub = 2.674402930e-18 lub = 5.724650092e-26   uc = 6.880685595e-11 luc = -5.441517696e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.565285543e-02 lu0 = -9.134878341e-10   a0 = 5.452179876e-01 la0 = 1.955396745e-7   keta = 2.186890623e-02 lketa = -9.878075601e-9   a1 = 0.0   a2 = 0.38689047   ags = 4.092176022e-01 lags = -8.253714428e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.318676412e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.082948430e-9   nfactor = {2.525307752e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.734922266e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.661000000e-07 lcit = 1.822092460e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.582008429e-03 leta0 = 5.788510789e-11   etab = 6.718111913e-03 letab = -3.090999436e-09 wetab = -9.305781891e-25 petab = 2.711709362e-31   dsub = 1.524923775e+00 ldsub = -2.371054445e-7   voffl = 0.0   minv = 0.0   pclm = 1.361199546e-01 lpclm = 8.524841786e-8   pdiblc1 = 0.39   pdiblc2 = 3.336387468e-03 lpdiblc2 = 1.810941255e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.876664321e-04 lalpha0 = 4.645703727e-10 walpha0 = 2.067951531e-25 palpha0 = -7.395570986e-32   alpha1 = 0.0   beta0 = 1.972811587e+01 lbeta0 = 2.058068375e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702362710e-01 lkt1 = -2.004301707e-10   kt2 = -4.492248858e-02 lkt2 = 4.121937564e-9   at = 1.041923757e+05 lat = -1.029700891e-2   ute = -1.217219698e+00 lute = 3.975805749e-8   ua1 = 1.721247906e-09 lua1 = -1.175978474e-16   ub1 = -1.641411537e-18 lub1 = 1.577822745e-25   uc1 = -2.697963625e-11 luc1 = 6.899025125e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.78 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.032128458e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.395290629e-07 wvth0 = -2.584759108e-07 pvth0 = 5.213329883e-14   k1 = -8.720072141e-02 lk1 = 1.387078140e-07 wk1 = 2.807599276e-07 pk1 = -5.662787360e-14   k2 = 5.372955957e-02 lk2 = -2.545693918e-08 wk2 = -5.448747510e-08 pk2 = 1.098985129e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.068828685e+05 lvsat = 7.620063618e-03 wvsat = 2.346971906e-02 pvsat = -4.733724985e-9   ua = 3.292517191e-09 lua = -1.105037891e-15 wua = -3.395211767e-15 pua = 6.847972374e-22   ub = 7.498483742e-18 lub = -9.157464785e-25 wub = -2.337536590e-24 pub = 4.714694425e-31   uc = -2.132339419e-10 luc = 5.144470103e-17 wuc = 1.745315453e-16 puc = -3.520214004e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.191608447e-01 lu0 = -1.977358174e-08 wu0 = -5.314109220e-08 pu0 = 1.071829259e-14   a0 = 4.364391664e+00 la0 = -5.747685602e-7   keta = 1.283487821e+00 lketa = -2.643403027e-07 wketa = -7.393984081e-07 pketa = 1.491329619e-13   a1 = 0.0   a2 = 0.38689047   ags = -2.003522107e+00 lags = 4.041003914e-07 wags = -3.521176466e-08 pags = 7.102036873e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-5.453977390e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.748990150e-08 wvoff = 2.464409033e-07 pvoff = -4.970589800e-14   nfactor = {-2.867426668e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.040338346e-06 wnfactor = 2.283039557e-06 pnfactor = -4.604776635e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 7.616524032e-05 lcit = -1.334519815e-11 wcit = -3.593037210e-11 pcit = 7.246976401e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.508009050e-01 leta0 = 3.099445184e-08 weta0 = 1.212565263e-08 peta0 = -2.445683507e-15   etab = -1.167955550e-01 letab = 2.182108961e-08 wetab = 8.203914313e-08 petab = -1.654688497e-14   dsub = 1.328602546e-01 ldsub = 4.366680724e-08 wdsub = 1.495091527e-07 pdsub = -3.015524856e-14   voffl = 0.0   minv = 0.0   pclm = 1.920727230e+00 lpclm = -2.746979465e-07 wpclm = -4.866409597e-07 ppclm = 9.815304838e-14   pdiblc1 = -1.166660283e+01 lpdiblc1 = 2.431756508e-06 wpdiblc1 = 6.905817518e-06 ppdiblc1 = -1.392868864e-12   pdiblc2 = -1.499775701e-02 lpdiblc2 = 5.508846525e-09 wpdiblc2 = 1.480331331e-08 ppdiblc2 = -2.985754277e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.557933004e-03 lalpha0 = -4.320848055e-10 walpha0 = -2.324287625e-10 palpha0 = 4.687971924e-17   alpha1 = 0.0   beta0 = 3.580275801e+01 lbeta0 = -1.184106570e-06 wbeta0 = -1.823574175e-06 pbeta0 = 3.678057933e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 1.894321030e-01 lkt1 = -9.291324286e-08 wkt1 = -2.523749336e-07 pkt1 = 5.090276224e-14   kt2 = -1.345778960e-01 lkt2 = 2.220498497e-08 wkt2 = 6.537171900e-08 pkt2 = -1.318514886e-14   at = -3.505321996e+04 lat = 1.778813150e-02 wat = 3.094323645e-02 pat = -6.241096077e-9   ute = 5.730355698e-01 lute = -3.213274788e-07 wute = -1.279121247e-07 pute = 2.579923599e-14   ua1 = 5.502381890e-09 lua1 = -8.802336663e-16 wua1 = -1.123039710e-15 pua1 = 2.265114944e-22   ub1 = -6.204888523e-18 lub1 = 1.078212765e-24 wub1 = 1.833311306e-24 pub1 = -3.697697239e-31   uc1 = -1.859700165e-10 luc1 = 3.896658986e-17 wuc1 = 1.181793055e-16 puc1 = -2.383617502e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.79 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-6.219809629e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.830887730e-08 wvth0 = 7.202888115e-07 pvth0 = -7.676512127e-14   k1 = 1.806557848e+00 lk1 = -1.106907209e-07 wk1 = -6.551064977e-07 pk1 = 6.662105529e-14   k2 = -3.619769999e-01 lk2 = 2.928953618e-08 wk2 = 1.300248201e-07 pk2 = -1.330949543e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.666708946e+05 lvsat = -2.537204751e-04 wvsat = 5.794577055e-03 pvsat = -2.405997159e-9   ua = -1.346939062e-08 lua = 1.102421559e-15 wua = 7.237541409e-15 pua = -7.154831921e-22   ub = -9.189124049e-18 lub = 1.281928030e-24 wub = 7.196493458e-24 pub = -7.841146447e-31   uc = 1.245358846e-09 luc = -1.406446761e-16 wuc = -7.130511725e-16 puc = 8.168806599e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.928823160e-01 lu0 = 2.132094231e-08 wu0 = 1.324068274e-07 pu0 = -1.371744069e-14   a0 = 0.0   keta = -2.962341822e+00 lketa = 2.948142322e-07 wketa = 1.724641454e-06 pketa = -1.753687677e-13   a1 = 0.0   a2 = 0.38689047   ags = 4.609831005e-01 lags = 7.953737810e-08 wags = 8.216078421e-08 pags = -8.355340950e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {8.021489523e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.997526000e-08 wvoff = -5.750417223e-07 pvoff = 5.847925639e-14   nfactor = {7.945692283e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.836953542e-07 wnfactor = -5.100504325e-06 pnfactor = 5.118981481e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.443855607e-04 lcit = 1.570023960e-11 wcit = 8.383753490e-11 pcit = -8.525858112e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.722625573e-01 leta0 = -2.472089084e-08 weta0 = -2.829318946e-08 peta0 = 2.877275903e-15   etab = 2.216874865e-01 letab = -2.275543454e-08 wetab = -1.914246673e-07 petab = 1.946693154e-14   dsub = 1.157306491e+00 ldsub = -9.124763988e-08 wdsub = -3.488546897e-07 pdsub = 3.547677767e-14   voffl = 0.0   minv = 0.0   pclm = -7.115775701e-01 lpclm = 7.196343410e-08 wpclm = 4.540484222e-07 ppclm = -2.573103978e-14   pdiblc1 = 2.645427494e+01 lpdiblc1 = -2.588572490e-06 wpdiblc1 = -1.611357421e-05 ppdiblc1 = 1.638669929e-12   pdiblc2 = -7.284274604e-02 lpdiblc2 = 1.312674236e-08 wpdiblc2 = 4.740609533e-08 ppdiblc2 = -7.279377656e-15   pdiblcb = 0.0   drout = 6.182016454e+01 ldrout = -7.681185222e-06 wdrout = -3.167311457e-05 pdrout = 4.171190823e-12   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.154137595e-03 lalpha0 = -1.155169692e-10 walpha0 = 5.705381554e-10 palpha0 = -5.886700901e-17   alpha1 = 0.0   beta0 = 2.830609109e+01 lbeta0 = -1.968330209e-07 wbeta0 = 1.788912857e-05 pbeta0 = -2.228258595e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -8.561658358e-01 lkt1 = 4.478677769e-08 wkt1 = 4.076044650e-07 pkt1 = -3.601322467e-14   kt2 = 2.154628732e-01 lkt2 = -2.389363414e-08 wkt2 = -1.525340110e-07 pkt2 = 1.551194625e-14   at = 2.206337314e+05 lat = -1.588456156e-02 wat = -1.098921762e-01 pat = 1.230622360e-8   ute = -2.351312646e+00 lute = 6.379455956e-08 wute = 2.984616243e-07 pute = -3.035205488e-14   ua1 = -6.647447783e-09 lua1 = 7.198381525e-16 wua1 = 4.032910689e-15 pua1 = -4.525013934e-22   ub1 = 7.521557381e-18 lub1 = -7.294915280e-25 wub1 = -4.277726381e-24 pub1 = 4.350233843e-31   uc1 = 4.180512706e-10 luc1 = -4.057999354e-17 wuc1 = -2.757517128e-16 puc1 = 2.804257043e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.80 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.741007788e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.737496073e-8   k1 = 7.034642523e-01 wk1 = -9.242771717e-8   k2 = -1.084412289e-01 wk2 = 2.781321683e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.465154812e+05 wvsat = -1.878730949e-1   ua = -3.168984913e-10 wua = -3.604040860e-16   ub = 1.024462025e-18 wub = 7.430622542e-25   uc = 1.332593942e-11 wuc = 4.900744622e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.558719343e-02 wu0 = 4.092320427e-9   a0 = 3.076023655e+00 wa0 = -6.262610184e-7   keta = 4.130400000e-01 wketa = -2.242972416e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.461445773e+00 wags = 2.156129010e-6   b0 = -3.063263502e-07 wb0 = 1.663474612e-13   b1 = -3.323065662e-09 wb1 = 1.804557577e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-4.693482038e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -3.437403538e-8   nfactor = {3.451418416e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.034756538e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.339746485e-01 weta0 = -1.379183931e-7   etab = -2.924061538e-01 wetab = 1.207754378e-7   dsub = 1.513169231e+00 wdsub = -5.176090191e-7   voffl = 0.0   minv = 0.0   pclm = 5.931222154e-02 wpclm = 7.639909122e-8   pdiblc1 = 0.39   pdiblc2 = -4.872617969e-03 wpdiblc2 = 6.756350526e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.065573686e-04 walpha0 = 8.052865361e-11   alpha1 = 0.0   beta0 = 4.742433271e+00 wbeta0 = 7.087176880e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.642704123e-01 wkt1 = 3.606009500e-9   kt2 = -5.101738831e-02 wkt2 = 7.957375987e-9   at = -2.695791138e+04 wat = 4.626044340e-2   ute = -1.576047508e+00 wute = 2.146352066e-7   ua1 = 1.504807877e-09 wua1 = 2.491424745e-16   ub1 = -9.820215385e-20 wub1 = -7.427689424e-25   uc1 = 1.447169809e-10 wuc1 = -4.414859860e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.81 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.741007788e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.737496073e-8   k1 = 7.034642523e-01 wk1 = -9.242771717e-8   k2 = -1.084412289e-01 wk2 = 2.781321683e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.465154812e+05 wvsat = -1.878730949e-1   ua = -3.168984913e-10 wua = -3.604040860e-16   ub = 1.024462025e-18 wub = 7.430622542e-25   uc = 1.332593942e-11 wuc = 4.900744622e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.558719343e-02 wu0 = 4.092320427e-9   a0 = 3.076023655e+00 wa0 = -6.262610184e-7   keta = 4.130400000e-01 wketa = -2.242972416e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.461445773e+00 wags = 2.156129010e-6   b0 = -3.063263502e-07 wb0 = 1.663474612e-13   b1 = -3.323065662e-09 wb1 = 1.804557577e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-4.693482038e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -3.437403538e-8   nfactor = {3.451418416e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.034756538e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.339746485e-01 weta0 = -1.379183931e-7   etab = -2.924061538e-01 wetab = 1.207754378e-7   dsub = 1.513169231e+00 wdsub = -5.176090191e-7   voffl = 0.0   minv = 0.0   pclm = 5.931222154e-02 wpclm = 7.639909122e-8   pdiblc1 = 0.39   pdiblc2 = -4.872617969e-03 wpdiblc2 = 6.756350526e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.065573686e-04 walpha0 = 8.052865361e-11   alpha1 = 0.0   beta0 = 4.742433271e+00 wbeta0 = 7.087176880e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.642704123e-01 wkt1 = 3.606009500e-9   kt2 = -5.101738831e-02 wkt2 = 7.957375987e-9   at = -2.695791138e+04 wat = 4.626044340e-2   ute = -1.576047508e+00 wute = 2.146352066e-7   ua1 = 1.504807877e-09 wua1 = 2.491424745e-16   ub1 = -9.820215385e-20 wub1 = -7.427689424e-25   uc1 = 1.447169809e-10 wuc1 = -4.414859860e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.82 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.437035099e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.201207355e-07 wvth0 = -1.481967278e-08 pvth0 = -4.961466859e-14   k1 = 1.010534960e+00 lk1 = -1.213449779e-06 wk1 = -2.192602022e-07 pk1 = 5.012032969e-13   k2 = -2.300874058e-01 lk2 = 4.807085892e-07 wk2 = 7.805795376e-08 pk2 = -1.985518757e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.189973935e+06 lvsat = -2.542751554e+00 wvsat = -4.536471747e-01 pvsat = 1.050258102e-6   ua = 2.189041438e-10 lua = -2.117328594e-15 wua = -5.817120064e-16 pua = 8.745414025e-22   ub = 2.625940407e-19 lub = 3.010669903e-24 wub = 1.057744206e-24 pub = -1.243527097e-30   uc = -1.053543128e-10 luc = 4.689881592e-16 wuc = 5.392043599e-17 puc = -1.937108693e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.466239413e-02 lu0 = 3.654524777e-09 wu0 = 4.474299530e-09 pu0 = -1.509464914e-15   a0 = 3.306481179e+00 la0 = -9.106978450e-07 wa0 = -7.214491941e-07 pa0 = 3.761546379e-13   keta = 1.151795135e+00 lketa = -2.919334973e-06 wketa = -5.294326626e-07 pketa = 1.205802117e-12   a1 = 0.0   a2 = 0.38689047   ags = -7.437045750e+00 lags = 1.571035855e-05 wags = 3.798210825e-06 pags = -6.489006496e-12   b0 = -3.063263502e-07 wb0 = 1.663474612e-13   b1 = -3.323065662e-09 wb1 = 1.804557577e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.919255338e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.096289778e-07 wvoff = -4.583270134e-08 pvoff = 4.528115298e-14   nfactor = {4.487451381e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.094086288e-06 wnfactor = -1.462679594e-06 pnfactor = 1.691021400e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 6.580436947e-01 leta0 = -1.280622029e-06 weta0 = -2.717718720e-07 peta0 = 5.289481230e-13   etab = -5.757117980e-01 letab = 1.119537497e-06 wetab = 2.377920010e-07 petab = -4.624137679e-13   dsub = 2.156240106e+00 ldsub = -2.541219963e-06 wdsub = -7.832230134e-07 pdsub = 1.049625493e-12   voffl = 0.0   minv = 0.0   pclm = -8.144380567e-02 lpclm = 5.562248890e-07 wpclm = 1.345369607e-07 ppclm = -2.297431281e-13   pdiblc1 = 0.39   pdiblc2 = -2.190723604e-02 lpdiblc2 = 6.731561507e-08 wpdiblc2 = 1.379232918e-08 ppdiblc2 = -2.780404165e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.436704710e-04 lalpha0 = 1.332168161e-09 walpha0 = 2.197698494e-10 palpha0 = -5.502387374e-16   alpha1 = 0.0   beta0 = -9.108448967e+00 lbeta0 = 5.473446209e-05 wbeta0 = 1.280814528e-05 pbeta0 = -2.260752222e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.198790675e-01 lkt1 = -1.754210553e-07 wkt1 = -1.472939156e-08 pkt1 = 7.245591270e-14   kt2 = -4.806204166e-02 lkt2 = -1.167862857e-08 wkt2 = 6.736699607e-09 pkt2 = 4.823740744e-15   at = 9.965578175e+03 lat = -1.459103691e-01 wat = 3.100956527e-02 pat = 6.026681884e-8   ute = -1.825111894e+00 lute = 9.842264904e-07 wute = 3.175087607e-07 pute = -4.065249096e-13   ua1 = 1.167694542e-09 lua1 = 1.332169080e-15 wua1 = 3.883837663e-16 pua1 = -5.502391166e-22   ub1 = 1.647694355e-18 lub1 = -6.899250505e-24 wub1 = -1.463894036e-24 pub1 = 2.849666429e-30   uc1 = 4.406922980e-10 luc1 = -1.169604181e-15 wuc1 = -1.663982436e-16 puc1 = 4.830933108e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.83 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.979705956e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.809615643e-07 wvth0 = -7.853814987e-08 pvth0 = 7.474436454e-14   k1 = 3.022876744e-01 lk1 = 1.688329063e-07 wk1 = 7.327425658e-08 pk1 = -6.973474362e-14   k2 = 7.076605000e-02 lk2 = -1.064655962e-07 wk2 = -4.620655763e-08 pk2 = 4.397454986e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3.075186907e+05 lvsat = 3.798973158e-01 wvsat = 1.648771795e-01 pvsat = -1.569127873e-7   ua = -5.580883861e-10 lua = -6.008761583e-16 wua = -2.607830118e-16 pua = 2.481858884e-22   ub = 8.360910974e-19 lub = 1.891378565e-24 wub = 8.208669819e-25 pub = -7.812150024e-31   uc = 2.393945250e-10 luc = -2.038564237e-16 wuc = -8.847462396e-17 puc = 8.420085725e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.800758206e-02 lu0 = 1.664268822e-08 wu0 = 7.223003108e-09 pu0 = -6.874095943e-15   a0 = 4.058091078e+00 la0 = -2.377611128e-06 wa0 = -1.031894147e-06 pa0 = 9.820485002e-13   keta = -5.476618172e-01 lketa = 3.974866631e-07 wketa = 1.725110370e-07 pketa = -1.641778913e-13   a1 = 0.0   a2 = 0.38689047   ags = -4.782324498e-01 lags = 2.128877428e-06 wags = 9.239425791e-07 pags = -8.793115328e-13   b0 = -6.896113760e-07 lb0 = 7.480554685e-13 wb0 = 3.246595083e-13 pb0 = -3.089768307e-19   b1 = -7.480988437e-09 lb1 = 8.114997091e-15 wb1 = 3.521946000e-15 pb1 = -3.351818398e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.321734584e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.017738104e-07 wvoff = -4.417030106e-08 pvoff = 4.203665466e-14   nfactor = {3.763558915e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.681268981e-06 wnfactor = -1.163683050e-06 pnfactor = 1.107471340e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.617510060e-03 leta0 = -3.381716906e-09 weta0 = -1.467680665e-09 peta0 = 1.396784351e-15   etab = -4.076340203e-03 letab = 3.879432590e-09 wetab = 1.683691557e-09 petab = -1.602360837e-15   dsub = 1.419662371e+00 ldsub = -1.103644880e-06 wdsub = -4.789869458e-07 pdsub = 4.558494814e-13   voffl = 0.0   minv = 0.0   pclm = 1.647913660e-01 lpclm = 7.564893550e-08 wpclm = 3.283198537e-08 ppclm = -3.124603632e-14   pdiblc1 = 0.39   pdiblc2 = 1.362915495e-02 lpdiblc2 = -2.040581542e-09 wpdiblc2 = -8.856217592e-10 ppdiblc2 = 8.428418002e-16   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.821209063e-04 lalpha0 = -2.795247409e-10 walpha0 = -1.213150211e-10 palpha0 = 1.154548990e-16   alpha1 = 0.0   beta0 = 1.611446988e+01 lbeta0 = 5.507017497e-06 wbeta0 = 2.390070881e-06 pbeta0 = -2.274618507e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.613617917e-01 lkt1 = 1.007100700e-07 wkt1 = 4.370863283e-08 pkt1 = -4.159728732e-14   kt2 = -7.526285533e-02 lkt2 = 4.140906346e-08 wkt2 = 1.797172368e-08 pkt2 = -1.710359957e-14   at = -2.073946462e+05 lat = 2.783104940e-01 wat = 1.207880323e-01 pat = -1.149533664e-7   ute = -1.572464670e+00 lute = 4.911361658e-07 wute = 2.131553512e-07 pute = -2.028588819e-13   ua1 = 1.604979619e-09 lua1 = 4.787219816e-16 wua1 = 2.077675382e-16 pua1 = -1.977313273e-22   ub1 = -1.878564103e-18 lub1 = -1.706950339e-26 wub1 = -7.408242853e-27 pub1 = 7.050387682e-33   uc1 = -3.455098480e-10 luc1 = 3.648226166e-16 wuc1 = 1.583346908e-16 puc1 = -1.506863336e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.84 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.927364836e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.435871391e-8   k1 = 4.858330520e-01 lk1 = -5.846311873e-9   k2 = -3.823938991e-02 lk2 = -2.725664082e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.086556317e+04 lvsat = 5.785871325e-2   ua = -5.973298911e-10 lua = -5.635302142e-16   ub = 2.843642699e-18 lub = -1.919825649e-26   uc = -3.328092712e-12 luc = 2.714147794e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.621327065e-02 lu0 = -1.020052459e-08 wu0 = -1.323488980e-23   a0 = 2.085283895e+00 la0 = -5.001003956e-7   keta = -2.474407000e-01 lketa = 1.117677270e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.142883192e+00 lags = -1.317320223e-6   b0 = 1.835115401e-07 lb0 = -8.289124509e-14   b1 = 1.990755601e-09 lb1 = -8.992143512e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.367772733e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.300604696e-9   nfactor = {-3.856568835e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.267518948e-06 pnfactor = 2.019483917e-28   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.451695000e-05 lcit = -4.298758730e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.326232148e-03 leta0 = 2.274912835e-09 weta0 = 3.877409121e-25 peta0 = -3.697785493e-32   etab = 1.129237500e-04 letab = -1.074689683e-10   dsub = -4.085086000e-01 ldsub = 6.362162921e-7   voffl = 0.0   minv = 0.0   pclm = 1.714938677e-01 lpclm = 6.927019818e-8   pdiblc1 = 0.39   pdiblc2 = 1.522449257e-02 lpdiblc2 = -3.558856378e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.104386292e-05 lalpha0 = 4.507657599e-11   alpha1 = 0.0   beta0 = 1.974783646e+01 lbeta0 = 2.049160683e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.418626754e-01 lkt1 = -1.301664144e-8   kt2 = -2.809778745e-02 lkt2 = -3.477695813e-9   at = 8.833575994e+04 lat = -3.134654866e-3   ute = -9.906332080e-01 lute = -6.258992711e-8   ua1 = 2.692583669e-09 lua1 = -5.563453549e-16   ub1 = -2.442508916e-18 lub1 = 5.196339553e-25   uc1 = 8.258032704e-11 luc1 = -4.258866249e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.85 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.924389336e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.067638425e-8   k1 = 3.699287364e-01 lk1 = 4.650708796e-8   k2 = -2.151299859e-02 lk2 = -1.028089141e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.704909201e+05 lvsat = -5.209362345e-3   ua = -1.569550012e-09 lua = -1.243832468e-16   ub = 2.674402930e-18 lub = 5.724650092e-26   uc = 6.880685595e-11 luc = -5.441517696e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.565285543e-02 lu0 = -9.134878341e-10   a0 = 5.452179876e-01 la0 = 1.955396745e-7   keta = 2.186890623e-02 lketa = -9.878075601e-9   a1 = 0.0   a2 = 0.38689047   ags = 4.092176022e-01 lags = -8.253714428e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.318676412e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.082948430e-9   nfactor = {2.525307752e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.734922266e-08 wnfactor = 8.470329473e-22   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.661000000e-07 lcit = 1.822092461e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.582008429e-03 leta0 = 5.788510789e-11   etab = 6.718111913e-03 letab = -3.090999436e-09 wetab = -7.237830360e-25 petab = 3.081487911e-31   dsub = 1.524923775e+00 ldsub = -2.371054445e-7   voffl = 0.0   minv = 0.0   pclm = 1.361199546e-01 lpclm = 8.524841786e-8   pdiblc1 = 0.39   pdiblc2 = 3.336387468e-03 lpdiblc2 = 1.810941255e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.876664321e-04 lalpha0 = 4.645703727e-10 walpha0 = 1.033975766e-25 palpha0 = -3.697785493e-32   alpha1 = 0.0   beta0 = 1.972811587e+01 lbeta0 = 2.058068375e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702362710e-01 lkt1 = -2.004301707e-10   kt2 = -4.492248858e-02 lkt2 = 4.121937564e-9   at = 1.041923757e+05 lat = -1.029700891e-2   ute = -1.217219698e+00 lute = 3.975805749e-8   ua1 = 1.721247906e-09 lua1 = -1.175978474e-16   ub1 = -1.641411537e-18 lub1 = 1.577822745e-25   uc1 = -2.697963625e-11 luc1 = 6.899025125e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.86 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.561489524e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.352637649e-8   k1 = 4.298144664e-01 lk1 = 3.442843564e-8   k2 = -4.660830708e-02 lk2 = -5.219293166e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.501020035e+05 lvsat = -1.097019811e-3   ua = -2.959714260e-09 lua = 1.560059313e-16   ub = 3.193945236e-18 lub = -4.754258461e-26   uc = 1.081632762e-10 luc = -1.337951089e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.130232198e-02 lu0 = -3.600699061e-11   a0 = 4.364391664e+00 la0 = -5.747685602e-7   keta = -7.810323655e-02 lketa = 1.028580574e-8   a1 = 0.0   a2 = 0.38689047   ags = -2.068364043e+00 lags = 4.171786856e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-9.158051863e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.042762755e-9   nfactor = {1.336756371e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.923756480e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.284716979e-01 leta0 = 2.649076241e-08 weta0 = 8.271806126e-24 peta0 = -2.366582716e-30   etab = 3.427829431e-02 letab = -8.649750424e-09 petab = 7.888609052e-31   dsub = 4.081791128e-01 ldsub = -1.186362986e-8   voffl = 0.0   minv = 0.0   pclm = 1.024585215e+00 lpclm = -9.395058284e-8   pdiblc1 = 1.050356357e+00 lpdiblc1 = -1.331905755e-7   pdiblc2 = 1.226232200e-02 lpdiblc2 = 1.062488921e-11   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.129918930e-03 lalpha0 = -3.457565069e-10   alpha1 = 0.0   beta0 = 3.244467357e+01 lbeta0 = -5.067977288e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.753125450e-01 lkt1 = 8.234289138e-10   kt2 = -1.419685779e-02 lkt2 = -2.075268539e-9   at = 2.192828500e+04 lat = 6.295246857e-3   ute = 3.374873143e-01 lute = -2.738185734e-7   ua1 = 3.434321139e-09 lua1 = -4.631161530e-16   ub1 = -2.828873301e-18 lub1 = 3.972873752e-25   uc1 = 3.165539877e-11 luc1 = -4.927368263e-18 wuc1 = 6.162975822e-33 puc1 = -7.346839693e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.87 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.41525e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.48e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.996598e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.996598e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {8.768522871e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -8.576140215e-08 wvth0 = -9.363759662e-08 pvth0 = 1.233160329e-14   k1 = 6.001890767e-01 lk1 = 1.199095135e-8   k2 = 1.338272101e-02 lk2 = -1.311981161e-08 wk2 = -7.381052276e-08 pk2 = 9.720476795e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.519236538e+05 lvsat = -1.336922051e-03 wvsat = 1.380291868e-02 pvsat = -1.817775375e-9   ua = -4.649984676e-10 lua = -1.725356650e-16 wua = 1.756362915e-16 pua = -2.313042141e-23   ub = 6.803608967e-18 lub = -5.229172496e-25 wub = -1.488200279e-24 pub = 1.959885357e-31   uc = -3.220931744e-10 luc = 4.328311238e-17 wuc = 1.381379725e-16 puc = -1.819208029e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 5.398978013e-02 lu0 = -4.340781791e-09 wu0 = -1.654595633e-09 pu0 = 2.179019719e-16   a0 = 0.0   keta = -5.225893273e-01 lketa = 6.882240146e-08 wketa = 3.997582592e-07 pketa = -5.264616394e-14   a1 = 0.0   a2 = 0.38689047   ags = 6.122809500e-01 lags = 6.415114329e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.567905055e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.771456647e-08 wvoff = 4.760837205e-12 pvoff = -6.269784557e-19   nfactor = {-7.221146112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.319408616e-06 wnfactor = 3.135695597e-06 pnfactor = -4.129554316e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.201610741e-01 leta0 = -1.942243050e-8   etab = -1.308181618e-01 letab = 1.309262737e-8   dsub = 5.148958220e-01 ldsub = -2.591768688e-8   voffl = 0.0   minv = 0.0   pclm = 1.245457767e-01 lpclm = 2.458011099e-8   pdiblc1 = -3.218629833e+00 lpdiblc1 = 4.290135609e-07 wpdiblc1 = 1.058791184e-22 ppdiblc1 = -3.786532345e-29   pdiblc2 = 1.445486617e-02 lpdiblc2 = -2.781222148e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.540906590e-03 lalpha0 = -3.998815268e-10 walpha0 = -7.255728793e-10 palpha0 = 9.555432034e-17   alpha1 = 0.0   beta0 = 1.406724442e+02 lbeta0 = -1.475985398e-05 wbeta0 = -4.313029582e-05 pbeta0 = 5.680044308e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.055683383e-01 lkt1 = -2.153103438e-8   kt2 = -6.542621600e-02 lkt2 = 4.671381791e-9   at = -9.404356855e+04 lat = 2.156816011e-02 wat = 6.099018473e-02 pat = -8.032102379e-9   ute = -1.801700050e+00 lute = 7.901706585e-9   ua1 = 1.954026797e-09 lua1 = -2.681687898e-16 wua1 = -6.380340672e-16 pua1 = 8.402589648e-23   ub1 = -3.558114700e-19 lub1 = 7.159749729e-26   uc1 = -8.974136490e-11 luc1 = 1.105997853e-17 wuc1 = -6.162975822e-33 puc1 = 7.346839693e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.281312791e-10   cgso = 2.281312791e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.202975e-11   cgdl = 2.202975e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.11821e-8   dwc = 3.48e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00106130856   mjs = 0.42197   pbs = 0.7477   cjsws = 2.834310656e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.575208208e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__nfet_01v8_lvt





















