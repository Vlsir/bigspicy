** Translated using xdm 2.6.0 on Nov_14_2022_16_05_18_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_MULT=1.052 SKY130_FD_PR__NFET_05V0_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_05V0_NVT__OVERLAP_MULT=1.3700 SKY130_FD_PR__NFET_05V0_NVT__AJUNCTION_MULT=1.3878e+0 
+ SKY130_FD_PR__NFET_05V0_NVT__PJUNCTION_MULT=1.2464e+0 SKY130_FD_PR__NFET_05V0_NVT__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__WINT_DIFF=3.2175e-8 SKY130_FD_PR__NFET_05V0_NVT__DLC_DIFF=-3.0000e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__DWC_DIFF=3.2175e-8 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_0=-0.056577 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_0=0.08428 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_0=0.00016793 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_0=-0.005636 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_0=-1.9616e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_0=0.032906 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_0=0.0068039 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_0=-1.0516e-18 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_1=-1.0828e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_1=0.091002 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_1=0.042279 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_1=-0.0025266 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_1=-0.0056151 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_1=-2.4885e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_1=0.020743 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_1=0.004878 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_2=-1.0026e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_2=-0.19806 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_2=0.0025007 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_2=-0.0058474 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_2=-1.9172e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_2=2871.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_2=0.040758 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_3=-1.2607e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_3=0.021014 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_3=-7.6708e-19 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_3=0.1208 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_3=0.00073216 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_3=-0.004008 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_3=-0.0057207 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_3=0.001698 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_4=-0.0061975 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_4=0.014978 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_4=-2.6745e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_4=0.033608 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_4=-1.0632e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_4=0.12546 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_4=0.1273 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_4=-0.001136 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_5=0.00076607 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_5=-0.0073364 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_5=0.012511 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_5=-1.8417e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_5=0.026896 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_5=-1.0258e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_5=0.12026 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_5=0.11694 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_6=0.062703 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_6=-0.0018694 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_6=-0.0057585 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_6=0.0066755 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_6=-1.5181e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_6=0.013027 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_6=-8.6079e-19 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_6=0.15139 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_7=-0.062415 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_7=0.00069645 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_7=-0.0070762 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_7=0.020702 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_7=-2.2827e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_7=3748.4 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_7=-1.0099e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_8=0.010794 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_8=-2.5551e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_8=0.0029018 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_8=-0.0068423 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_8=0.0021841 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_8=-6.2851e-12 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_8=3.5554e-10 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_8=-6.4524e-19 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_9=0.15402 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_9=0.004958 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_9=-0.0072966 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_9=0.035399 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_9=2.2764e-13 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_9=1592.8 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_9=-2.896e-19 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_10=2509.5 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_10=0.025399 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_10=-0.019006 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_10=-0.0078678 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_10=0.00080055 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_10=-1.5105e-11 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_10=-7.9876e-19 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0, L = 2.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0, L = 4.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0, L = 0.9
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0, L = 25.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0, L = 2.0
* ------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0, L = 4.0
* ------------------------------------
*














* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0, L = 8.0
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0, L = 0.9
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42, L = 1.0
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42, L = 0.9
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7, L = 0.9
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_05v0_nvt.pm3.spice




















