** Translated using xdm 2.6.0 on Nov_14_2022_16_05_32_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__RF_PFET_01V8_B__TOXE_MULT=1.052 SKY130_FD_PR__RF_PFET_01V8_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_PFET_01V8_B__OVERLAP_MULT=1.1934 SKY130_FD_PR__RF_PFET_01V8_B__AJUNCTION_MULT=1.0909 
+ SKY130_FD_PR__RF_PFET_01V8_B__PJUNCTION_MULT=1.096 SKY130_FD_PR__RF_PFET_01V8_B__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__RF_PFET_01V8_B__WINT_DIFF=3.2175e-8 SKY130_FD_PR__RF_PFET_01V8_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__DLC_DIFF=-1.7325e-8 SKY130_FD_PR__RF_PFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__XGW_DIFF=6.4250e-8 SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT=1.15 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT=1.45 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT=1.45 
+ SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT_2=1.15 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT_2=1.30 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT_2=1.30 SKY130_FD_PR__RF_PFET_01V8__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RS_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_0=-0.026318 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_0=-0.00026051 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_0=0.036371 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_0=9011.9 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_1=-0.0083086 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_1=-0.00025544 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_1=0.043744 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_1=-13691.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_2=0.00092097 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_2=-0.00036227 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_2=0.025821 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_2=-12946.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_3=-0.023482 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_3=-0.00065054 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_3=0.062883 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_3=-10906.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_4=-0.018913 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_4=-0.00048132 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_4=0.054592 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_4=-4787.1 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_5=-0.016498 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_5=-0.00040228 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_5=0.025581 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_5=-7701.6 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_6=-0.02415 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_6=-0.0010764 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_6=0.088259 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_6=-9692.8 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_7=-0.00045958 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_7=-12867.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_7=-0.013677 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_7=0.054734 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_8=0.03218 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_8=-0.00053308 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_8=-16884.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_8=-0.012368 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_0=-0.025153 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_0=-0.00045786 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_0=0.049883 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_0=4304.4 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_1=-0.0081868 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_1=-0.0003546 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_1=0.058034 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_1=-1647.5 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_2=-0.00039936 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_2=0.0326 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_2=-10830.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_2=-0.00049705 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_3=-0.021287 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_3=-0.00070687 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_3=0.061799 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_3=-10201.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_4=-0.00073938 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_4=0.067454 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_4=-10506.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_4=-0.015399 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_5=0.033162 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_5=-0.00052171 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_5=-14143.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_5=-0.016662 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_6=0.091648 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_6=-0.00096119 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_6=-7280.9 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_6=-0.023369 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_7=-0.010709 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_7=0.059069 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_7=-0.0007366 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_7=-12730.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_8=-0.0113 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_8=0.044518 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_8=-0.00066793 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_8=-13679.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_8=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_pfet_01v8_b.pm3.spice














