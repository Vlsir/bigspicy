** Translated using xdm 2.6.0 on Nov_14_2022_16_05_12_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
.PARAM 
+ SKY130_FD_PR__NFET_01V8_LVT__LKVTH0_DIFF=0.0 SKY130_FD_PR__NFET_01V8_LVT__WLOD_DIFF=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__LKU0_DIFF=0.0 SKY130_FD_PR__NFET_01V8_LVT__KVTH0_DIFF=7.9e-9 
+ SKY130_FD_PR__NFET_01V8_LVT__WKVTH0_DIFF=.3e-6 SKY130_FD_PR__NFET_01V8_LVT__KU0_DIFF=-2.7e-8 
+ SKY130_FD_PR__NFET_01V8_LVT__WKU0_DIFF=0.0 SKY130_FD_PR__NFET_01V8_LVT__KVSAT_DIFF=0.2 
+ SKY130_FD_PR__PFET_01V8__LKVTH0_DIFF=.0e-6 SKY130_FD_PR__PFET_01V8__WLOD_DIFF=.0e-6 
+ SKY130_FD_PR__PFET_01V8__LKU0_DIFF=0.0 SKY130_FD_PR__PFET_01V8__KVSAT_DIFF=0.5 
+ SKY130_FD_PR__PFET_01V8__KVTH0_DIFF=3.29e-8 SKY130_FD_PR__PFET_01V8__WKVTH0_DIFF=.20e-6 
+ SKY130_FD_PR__PFET_01V8__KU0_DIFF=4.5e-8 SKY130_FD_PR__PFET_01V8__WKU0_DIFF=.25e-6 
+ SKY130_FD_PR__PFET_01V8_LVT__WKVTH0_DIFF=.73e-6 SKY130_FD_PR__PFET_01V8_LVT__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__WLOD_DIFF=.0e-6 SKY130_FD_PR__PFET_01V8_LVT__KU0_DIFF=5.9e-8 
+ SKY130_FD_PR__PFET_01V8_LVT__LKU0_DIFF=0.0 SKY130_FD_PR__PFET_01V8_LVT__WKU0_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KVSAT_DIFF=.0e-6 SKY130_FD_PR__PFET_01V8_LVT__KVTH0_DIFF=1.76e-8 
+ SKY130_FD_PR__NFET_G5V0D10V5__WKVTH0_DIFF=.65e-6 SKY130_FD_PR__NFET_G5V0D10V5__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KVTH0_DIFF=11.0e-9 SKY130_FD_PR__NFET_G5V0D10V5__WLOD_DIFF=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KU0_DIFF=-4.5e-8 SKY130_FD_PR__NFET_G5V0D10V5__LKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__WKU0_DIFF=.2e-6 SKY130_FD_PR__NFET_G5V0D10V5__KVSAT_DIFF=0.3 
+ SKY130_FD_PR__PFET_G5V0D10V5__WKVTH0_DIFF=.65e-6 SKY130_FD_PR__PFET_G5V0D10V5__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KVTH0_DIFF=3.5e-8 SKY130_FD_PR__PFET_G5V0D10V5__WLOD_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KU0_DIFF=7.0e-8 SKY130_FD_PR__PFET_G5V0D10V5__LKU0_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__WKU0_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KVSAT_DIFF=0.4 
+ SKY130_FD_PR__NFET_05V0_NVT__WKVTH0_DIFF=.8e-6 SKY130_FD_PR__NFET_05V0_NVT__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KVTH0_DIFF=-7.0e-9 SKY130_FD_PR__NFET_05V0_NVT__WLOD_DIFF=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KU0_DIFF=-3.0e-8 SKY130_FD_PR__NFET_05V0_NVT__LKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__WKU0_DIFF=.2e-6 SKY130_FD_PR__NFET_05V0_NVT__KVSAT_DIFF=0.4 
+ SKY130_FD_PR__NFET_03V3_NVT__WKVTH0_DIFF=.0e-6 SKY130_FD_PR__NFET_03V3_NVT__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KVTH0_DIFF=-2.0e-9 SKY130_FD_PR__NFET_03V3_NVT__WLOD_DIFF=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KU0_DIFF=-3.0e-8 SKY130_FD_PR__NFET_03V3_NVT__LKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__WKU0_DIFF=.5e-6 SKY130_FD_PR__NFET_03V3_NVT__KVSAT_DIFF=0.3
.PARAM 
+ SKY130_FD_PR__NFET_G5V0D16V0__WKU0_DIFF=.2e-6 SKY130_FD_PR__NFET_G5V0D16V0__KVSAT_DIFF=0.3 
+ SKY130_FD_PR__NFET_G5V0D16V0__KVTH0_DIFF=1.7057e-8 SKY130_FD_PR__NFET_G5V0D16V0__KU0_DIFF=-9.9000e-8 
+ SKY130_FD_PR__NFET_G5V0D16V0__LKU0_DIFF=9.6975e-7 SKY130_FD_PR__NFET_G5V0D16V0__LKVTH0_DIFF=2.2691e-7 
+ SKY130_FD_PR__NFET_G5V0D16V0__WKVTH0_DIFF=2.3093e-6
























* parameters fixed copy from Hvnmos
* parameters fixed copy from Hvpmos







.PARAM 
+ SKY130_FD_PR__PFET_G5V0D16V0__WKU0_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D16V0__KVSAT_DIFF=0.4 
+ SKY130_FD_PR__PFET_G5V0D16V0__KVTH0_DIFF=5.2302e-9 SKY130_FD_PR__PFET_G5V0D16V0__KU0_DIFF=2.2180e-7 
+ SKY130_FD_PR__PFET_G5V0D16V0__LKU0_DIFF=8.7129e-7 SKY130_FD_PR__PFET_G5V0D16V0__LKVTH0_DIFF=-4.8631e-7 
+ SKY130_FD_PR__PFET_G5V0D16V0__WKVTH0_DIFF=5.3980e-7
