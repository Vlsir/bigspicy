** Translated using xdm 2.6.0 on Nov_14_2022_16_05_33_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

*
* model corner
* , Bin 000, W = 30.0, L = 1.0
* ----------------------------
.PARAM 
+ SKY130_FD_PR__NFET_20V0_NVT__RDRIFT_MULT=7.2610e-1 SKY130_FD_PR__NFET_20V0_NVT__HVVSAT_MULT=5.4501e-1 
+ SKY130_FD_PR__NFET_20V0_NVT__VTH0_DIFF=3.0654e-2 SKY130_FD_PR__NFET_20V0_NVT__K2_DIFF=-1.2365e-1
.INCLUDE sky130_fd_pr__nfet_20v0_nvt__subcircuit.pm3.spice


