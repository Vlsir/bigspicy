** Translated using xdm 2.6.0 on Nov_14_2022_16_05_02_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM 
+ SKY130_FD_PR__NFET_20V0__TOXE_MULT=1.06 SKY130_FD_PR__NFET_20V0__RSHN_MULT=1.0 SKY130_FD_PR__NFET_20V0__OVERLAP_MULT=0.10 
+ SKY130_FD_PR__NFET_20V0__AJUNCTION_MULT=1.6 SKY130_FD_PR__NFET_20V0__PJUNCTION_MULT=1.6 
+ SKY130_FD_PR__NFET_20V0__LINT_DIFF=-1.7325e-8 SKY130_FD_PR__NFET_20V0__WINT_DIFF=3.2175e-8 
+ SKY130_FD_PR__NFET_20V0__DLC_DIFF=-1.7325e-8 SKY130_FD_PR__NFET_20V0__DWC_DIFF=3.2175e-8
.PARAM 
+ SKY130_FD_PR__NFET_20V0__RDRIFT_MULT=1.8205 SKY130_FD_PR__NFET_20V0__HVVSAT_MULT=1.3172 
+ SKY130_FD_PR__NFET_20V0__VTH0_DIFF=1.7977e-1 SKY130_FD_PR__NFET_20V0__K2_DIFF=-2.5783e-2



.PARAM 
+ SKY130_FD_PR__NFET_20V0_ISO__RDRIFT_MULT=2.3846 SKY130_FD_PR__NFET_20V0_ISO__HVVSAT_MULT=2.4860 
+ SKY130_FD_PR__NFET_20V0_ISO__VTH0_DIFF=1.4387e-1 SKY130_FD_PR__NFET_20V0_ISO__K2_DIFF=-1.9447e-2


.INCLUDE sky130_fd_pr__nfet_20v0__subcircuit.pm3.spice




.INCLUDE sky130_fd_pr__nfet_20v0_iso__subcircuit.pm3.spice
.INCLUDE sky130_fd_pr__nfet_20v0_zvt__fs_discrete.corner.spice
