** Translated using xdm 2.6.0 on Nov_14_2022_16_05_34_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 2
.PARAM 
+ SKY130_FD_PR__PFET_01V8_MVT__TOXE_MULT=1.0 SKY130_FD_PR__PFET_01V8_MVT__RSHP_MULT=1.0 
+ SKY130_FD_PR__PFET_01V8_MVT__OVERLAP_MULT=9.5435e-1 SKY130_FD_PR__PFET_01V8_MVT__AJUNCTION_MULT=9.9626e-1 
+ SKY130_FD_PR__PFET_01V8_MVT__PJUNCTION_MULT=1.0009 SKY130_FD_PR__PFET_01V8_MVT__WINT_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__LINT_DIFF=0.0 SKY130_FD_PR__PFET_01V8_MVT__DLC_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__DWC_DIFF=0.0 SKY130_FD_PR__RF_PFET_01V8_MVT__AW_CAP_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RGATE_DIST_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RGATE_STUB_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RGATE_DIST_MULT_2=1.0 SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RGATE_STUB_MULT_2=1.0 
+ SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RD_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RS_MULT=1.0 
+ SKY130_FD_PR__PFET_01V8_MVT__B0_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__PDITSD_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__UA_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__U0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__B1_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__AGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__UB_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__KETA_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__K2_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__VTH0_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__A0_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__A0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__B0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__UA_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__U0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__TVOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__B1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__AGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__UB_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__K2_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__VTH0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__NFACTOR_DIFF_1=0.0
*
* sky130_fd_pr__pfet_01v8_mvt, Bin 000, W = 1.68, L = 0.15
* ------------------------------------
*








* sky130_fd_pr__pfet_01v8_mvt, Bin 001, W = 0.84, L = 0.15
* ------------------------------------
.INCLUDE sky130_fd_pr__pfet_01v8_mvt.pm3.spice























