** Translated using xdm 2.6.0 on Nov_14_2022_16_05_20_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_B__TOXE_MULT=0.9635 SKY130_FD_PR__RF_NFET_01V8_B__RBPB_MULT=0.8 
+ SKY130_FD_PR__RF_NFET_01V8_B__OVERLAP_MULT=0.95013 SKY130_FD_PR__RF_NFET_01V8_B__AJUNCTION_MULT=8.4039e-1 
+ SKY130_FD_PR__RF_NFET_01V8_B__PJUNCTION_MULT=8.6147e-1 SKY130_FD_PR__RF_NFET_01V8_B__LINT_DIFF=1.21275e-8 
+ SKY130_FD_PR__RF_NFET_01V8_B__WINT_DIFF=-2.252e-8 SKY130_FD_PR__RF_NFET_01V8_B__RSHG_DIFF=-7.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__DLC_DIFF=8.0874e-9 SKY130_FD_PR__RF_NFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__XGW_DIFF=-4.504e-8 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_0=-0.056554 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_0=-10484.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_0=0.0088666 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_0=0.0032864 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_1=-0.026928 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_1=-10520.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_1=0.019351 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_1=0.0032695 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_2=-0.032372 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_2=-8970.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_2=0.036836 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_2=0.0021845 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_3=-0.021269 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_3=-18297.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_3=0.008336 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_3=-0.001876 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_4=-0.040313 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_4=-16962.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_4=0.02702 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_4=-0.0017137 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_5=-0.024547 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_5=-13923.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_5=0.041021 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_5=0.0023309 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_6=-0.0015646 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_6=-0.029946 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_6=-19400.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_6=0.0046177 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_7=0.023534 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_7=-0.0020753 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_7=-0.036064 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_7=-15473.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_8=0.039622 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_8=9.7301e-5 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_8=-0.02617 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_8=-10255.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_0=0.0079125 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_0=0.0019161 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_0=-0.032091 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_0=-19913.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_1=0.02665 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_1=0.00077838 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_1=-0.04404 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_1=-14015.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_2=0.040538 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_2=0.001113 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_2=-0.035283 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_2=-10762.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_3=-20443.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_3=0.010632 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_3=-0.0029861 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_3=-0.031657 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_4=-16322.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_4=0.031114 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_4=-0.0056646 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_4=-0.048693 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_5=-950.61 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_5=0.043251 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_5=-0.0032668 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_5=-0.032962 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_6=-20376.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_6=0.006878 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_6=-0.0015387 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_6=-0.032585 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_7=-0.0046032 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_7=-19465.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_7=0.028329 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_7=-0.049601 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_8=-0.031697 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_8=-0.0020892 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_8=-5015.2 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_8=0.041815
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*





* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_b.pm3.spice














