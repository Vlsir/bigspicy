** Translated using xdm 2.6.0 on Nov_14_2022_16_05_05_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PFET_01V8__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__pfet_01v8 d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__pfet_01v8 d g s b sky130_fd_pr__pfet_01v8__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__pfet_01v8__model.0 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.069709+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43448553   k2 = 0.017927346   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.6228131e-10   ub = 1.00718446e-18   uc = -6.6549964e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0106298   a0 = 1.34499   keta = 0.0051290095   a1 = 0.0   a2 = 0.9995   ags = 0.1373328   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.23556545+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.3238158+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0015228006   pdiblc1 = 0.39   pdiblc2 = 0.0029632464   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.3760948e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.6464006   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1181082000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4485   kt2 = -0.0075706   at = 90900.0   ute = -0.33954   ua1 = 1.6104e-9   ub1 = -5.609e-19   uc1 = -1.0858e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.1 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.069709+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43448553   k2 = 0.017927346   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.6228131e-10   ub = 1.00718446e-18   uc = -6.6549964e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0106298   a0 = 1.34499   keta = 0.0051290095   a1 = 0.0   a2 = 0.9995   ags = 0.1373328   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.23556545+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.3238158+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0015228006   pdiblc1 = 0.39   pdiblc2 = 0.0029632464   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.3760948e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.6464006   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1181082000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4485   kt2 = -0.0075706   at = 90900.0   ute = -0.33954   ua1 = 1.6104e-9   ub1 = -5.609e-19   uc1 = -1.0858e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.2 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.07256076601125+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.29631129017263e-8   k1 = 0.438155474264772 lk1 = -2.95512830164046e-8   k2 = 0.016420547806151 lk2 = 1.21331052088333e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 268583.36765625 lvsat = -0.871823336188966   ua = -5.73170102295907e-10 lua = 8.76792015431752e-17   ub = 1.02351022777387e-18 lub = -1.31459049276751e-25   uc = -7.3265596390909e-11 luc = 5.40759039102703e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01053518012595 lu0 = 7.61902218480005e-10   a0 = 1.47724609397325 la0 = -1.06495820690344e-6   keta = 0.0215551457611434 lketa = -1.32267240725838e-07 wketa = 1.32348898008484e-23   a1 = 0.0   a2 = 1.201605619625 la2 = -1.62740356088607e-6   ags = 0.0295086516120699 lags = 8.68226244087671e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.242968604173382+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.96119963705402e-8   nfactor = {1.15676988289277+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.34509431670523e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.436220819781416 lpclm = 3.52481800301092e-06 wpclm = 1.32348898008484e-22 ppclm = -8.45658890396925e-28   pdiblc1 = 0.39   pdiblc2 = 0.00580619790136215 lpdiblc2 = -2.28921363261828e-8   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.01463321822624e-08 lpscbe2 = -6.20213856966074e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.23603180931265 lbeta0 = 1.13566322222307e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 8.41723541969075e-11 lagidl = 1.27448050124431e-16   bgidl = 1364529066.7315 lbgidl = -1477.16035895925   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.431471725249045 lkt1 = -1.37115806165454e-7   kt2 = 0.00990843714472826 lkt2 = -1.40745454495378e-7   at = 87841.8025997225 lat = 0.0246253486090028   ute = -0.47523588096623 lute = 1.09265620763916e-6   ua1 = 1.22154240555877e-09 lua1 = 3.13117584283619e-15   ub1 = -2.9782157667176e-19 lub1 = -2.11837139269586e-24   uc1 = -8.818088717071e-11 luc1 = -1.64258613485861e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.3 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.07437596491725+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.03187399621725e-8   k1 = 0.424193366780375 lk1 = 2.70265693024933e-8   k2 = 0.021758652454319 lk2 = -9.49819198497299e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53437.5   ua = -2.24827727670615e-10 lua = -1.32388874763554e-15   ub = 7.81807564174605e-19 lub = 8.47978877374716e-25   uc = -8.1142522719913e-11 luc = 8.59951234884924e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0121388372214 lu0 = -5.7365060209576e-9   a0 = 1.228324476138 la0 = -5.62673234818787e-8   keta = -0.005397538898584 lketa = -2.30484129822503e-8   a1 = 0.0   a2 = 0.8   ags = 0.0529089695462651 lags = 7.73402469541054e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.235249824251935+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.8333624465314e-8   nfactor = {1.4833449733681+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.17326923522308e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.16157665925 leta0 = -3.30568446409198e-7   etab = -0.141315443808768 letab = 2.88987507965972e-7   dsub = 0.86783645 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = 0.464982589871315 lpclm = -1.27077205330497e-7   pdiblc1 = 0.39   pdiblc2 = -2.37240050092149e-05 lpdiblc2 = 7.32123909457167e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800451626.855795 lpscbe1 = -1.83010176500738   pscbe2 = 8.28249481999155e-09 lpscbe2 = 1.35058333473979e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.8693587765981 lbeta0 = 8.79023745233698e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.31655291606185e-10 lagidl = -6.49643506117519e-17   bgidl = 916262739.3196 lbgidl = 339.323728431326   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.466380103196935 lkt1 = 4.34142401523773e-9   kt2 = -0.00524693839780851 lkt2 = -7.93321900407623e-8   at = 107195.154781301 lat = -0.0537991372953335   ute = -0.175352702489855 lute = -1.22543303159482e-7   ua1 = 2.34944805762225e-09 lua1 = -1.43937194039846e-15   ub1 = -1.03403519912063e-18 lub1 = 8.64945105377219e-25   uc1 = -2.43879612721223e-10 luc1 = 4.66670457235129e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.4 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0794830531205+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.07997259776741e-8   k1 = 0.35258842964425 lk1 = 1.73977300305546e-7   k2 = 0.050249560513596 lk2 = -6.79684586132678e-08 pk2 = 5.04870979341448e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 34694.4215625 lvsat = 0.0384653515218103   ua = -7.4590754973592e-10 lua = -2.54506330360777e-16   ub = 1.17217966544588e-18 lub = 4.68404651454509e-26   uc = -4.3075487117715e-11 luc = 7.87231614313079e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0101597196708 lu0 = -1.67487588156161e-9   a0 = 1.351594511058 la0 = -3.09247389756203e-7   keta = -0.006446117064797 lketa = -2.08964757806868e-8   a1 = 0.0   a2 = 0.6947757 la2 = 2.159458331049e-7   ags = 0.30333918616215 lags = 2.59458810502621e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.2342745959177+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.63322189429783e-8   nfactor = {1.2668641330019+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.66003981627882e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.5145729485 leta0 = 1.05705485304849e-06 weta0 = 2.13412598038681e-22 peta0 = 1.57772181044202e-28   etab = 7.82572104062834 letab = -1.60613073479647e-05 wetab = 1.22091858412827e-21 petab = 1.18944447289224e-26   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = 0.17740276109201 lpclm = 4.6310648522303e-7   pdiblc1 = 0.40904087372893 lpdiblc1 = -3.90764998240805e-8   pdiblc2 = 0.00023097199624504 lpdiblc2 = 2.0942582375513e-10   pdiblcb = -0.0505225220816911 lpdiblcb = 5.23784172844961e-8   drout = 0.39628460522442 ldrout = 3.35983772920421e-7   pscbe1 = 799096746.28841 lpscbe1 = 0.950442395244636   pscbe2 = 8.9459351914306e-09 lpscbe2 = -1.09575234634111e-17   pvag = 0.0   delta = 0.01   alpha0 = -4.6979642602591e-05 lalpha0 = 9.64138478979692e-11 walpha0 = -1.74882574078446e-26 palpha0 = -3.49601423889355e-33   alpha1 = 2.052243e-10 lalpha1 = -2.159458331049e-16   beta0 = -14.725699412172 lbeta0 = 4.69518154548331e-05 pbeta0 = 2.58493941422821e-26   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 791118977.9994 lbgidl = 596.149136594378   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.45601487547626 lkt1 = -1.69305420179237e-8   kt2 = -0.040265285984791 lkt2 = -7.46603133381056e-9   at = 70618.830790588 lat = 0.0212643675803393   ute = -0.16301041967218 lute = -1.47872666676076e-7   ua1 = 1.4104394005622e-09 lua1 = 4.87702002992429e-16   ub1 = 5.28204025400006e-21 lub1 = -1.26798642390869e-24   uc1 = -2.1727509487971e-11 luc1 = 1.07603584394091e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.5 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0794679540578+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.07838380946417e-8   k1 = 0.56491536311668 lk1 = -4.94422291522848e-8   k2 = -0.036353830017708 lk2 = 2.31593528495631e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 75015.192774 lvsat = -0.00396189774009209   ua = -6.571121372545e-10 lua = -3.47940681576463e-16   ub = 1.12564882108724e-18 lub = 9.58022204059194e-26   uc = -6.0433515316068e-11 luc = 2.61371798086503e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0102728845896 lu0 = -1.79395287521447e-9   a0 = 1.220834686686 la0 = -1.71656279879537e-7   keta = -0.04409425524965 lketa = 1.87185140873575e-08 wketa = -5.29395592033938e-23   a1 = 0.0   a2 = 1.0104486 la2 = -1.162187662098e-7   ags = 0.23070757605774 lags = 3.35884913813716e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17620407007814+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.47720853780177e-8   nfactor = {2.4585388898312+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.87927439522452e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -15.6534252956466 letab = 8.64446003035627e-6   dsub = 0.21654111562154 ldsub = 4.57293068750438e-8   voffl = 0.0   minv = 0.0   pclm = 0.61134393685442 lpclm = 6.49492061526446e-9   pdiblc1 = 0.739755433239658 lpdiblc1 = -3.87068580067328e-7   pdiblc2 = 0.00043   pdiblcb = 0.246942244163382 lpdiblcb = -2.60626800743519e-07 wpdiblcb = -3.30872245021211e-23 ppdiblcb = 1.49094711086771e-28   drout = 0.40145694955116 ldrout = 3.30541209809019e-7   pscbe1 = 800000000.0   pscbe2 = 8.7029855369806e-09 lpscbe2 = 2.44684549784024e-16   pvag = 0.0   delta = 0.01   alpha0 = 9.3959585205182e-05 lalpha0 = -5.18884679881653e-11   alpha1 = -1.104486e-10 lalpha1 = 1.162187662098e-16   beta0 = 52.5267536657712 lbeta0 = -2.38141075292611e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1734776774.4006 lbgidl = -396.808174064211   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.43195105370738 lkt1 = -4.22515300274755e-8   kt2 = -0.03871541994061 lkt2 = -9.09686702973771e-9   at = 108308.62589584 lat = -0.0183944554905964   ute = -0.22986253790638 lute = -7.7527993228967e-8   ua1 = 3.4411459828964e-09 lua1 = -1.64909478332266e-15   ub1 = -2.9809874963314e-18 lub1 = 1.87429479207654e-24 pub1 = 1.40129846432482e-45   uc1 = -5.1065622173484e-11 luc1 = 4.16311821459513e-17 wuc1 = -2.46519032881566e-32 puc1 = -2.35098870164458e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.6 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0226664694244+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 9.41561581623903e-9   k1 = 0.0532166322842398 lk1 = 2.33139813058815e-7   k2 = 0.15099510310196 lk2 = -8.03027840232417e-08 wk2 = 6.61744490042422e-23 pk2 = 3.15544362088405e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 66665.879216 lvsat = 0.000648952227118513   ua = -4.258654214796e-10 lua = -4.75645061636141e-16   ub = 4.573918093368e-19 lub = 4.64842477346018e-25   uc = -2.90636747570015e-11 luc = 8.81340494878976e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0097443452056 lu0 = -1.50207070017616e-9   a0 = 1.21778863919204 la0 = -1.6997412147333e-7   keta = 0.076539893930312 lketa = -4.79008503582323e-08 pketa = 6.31088724176809e-30   a1 = 0.0   a2 = 0.8   ags = -0.623380510596121 lags = 8.07549081051703e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.25841574363812+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.06287358637663e-8   nfactor = {-0.623740948461601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 9.1424002521588e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.0803678193867 leta0 = -3.26026495681568e-7   etab = 0.0059473210899072 letab = -3.31888162815362e-09 wetab = -6.20385459414771e-25 petab = -2.46519032881566e-31   dsub = 0.1575810144388 ldsub = 7.82896100325038e-8   voffl = 0.0   minv = 0.0   pclm = 0.44235608619416 lpclm = 9.98172782274386e-8   pdiblc1 = -0.424734191462636 lpdiblc1 = 2.56012663747142e-07 ppdiblc1 = -1.76704842769507e-28   pdiblc2 = -0.011249839804896 lpdiblc2 = 6.45010977337518e-09 wpdiblc2 = -4.96308367531817e-24 ppdiblc2 = -1.18329135783152e-30   pdiblcb = -0.4063458 lpdiblcb = 1.001469486294e-7   drout = 1.64219348607812 ldrout = -3.54646857332239e-7   pscbe1 = 800004279.76088 lpscbe1 = -0.00236346798760678   pscbe2 = 9.46592034447e-09 lpscbe2 = -1.76640857108347e-16   pvag = 0.0   delta = 0.01   alpha0 = -9.61787712479e-09 lalpha0 = 5.36662961702541e-15 walpha0 = -3.94430452610506e-31 palpha0 = -1.59867231711831e-36   alpha1 = 2.208972e-10 lalpha1 = -6.67646324196e-17   beta0 = 1.92328807828559 lbeta0 = 4.13130211716873e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 355970457.3032 lbgidl = 364.627962908609   cgidl = 582.916182590424 lcgidl = -0.000156238481422284   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.44747945232 lkt1 = -3.36760805924462e-8   kt2 = 0.025537478384 lkt2 = -4.45800803592153e-8   at = 60492.336 lat = 0.008011755890352   ute = -0.379015047 lute = 4.84043585042105e-9   ua1 = 8.422641802e-10 lua1 = -2.13880499956189e-16   ub1 = 4.3749795216e-19 lub1 = -1.35398674546949e-26   uc1 = 7.79939761999999e-12 luc1 = 9.12338702013834e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.7 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.9762324106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.61875342502448e-9   k1 = 0.168957125018572 lk1 = 1.98158059313312e-7   k2 = 0.127825573179914 lk2 = -7.32999557910128e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 50605.8123514286 lvsat = 0.00550299501646717   ua = -1.16568444868571e-09 lua = -2.52039939396284e-16   ub = 1.24185936780857e-18 lub = 2.27742649070834e-25   uc = -9.86218093027713e-14 luc = 5.89204507184635e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00690456690814286 lu0 = -6.43767588217822e-10   a0 = 1.06642640588557 la0 = -1.24225945992083e-7   keta = -0.276257369333443 lketa = 5.87296528823947e-8   a1 = 0.0   a2 = 0.893879952843286 la2 = -2.83745585872132e-8   ags = 4.69761336268 lags = -8.00684070188891e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.057333193323286+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.01470573910401e-8   nfactor = {4.11868964855714+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -5.19126425718857e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.559502569681777 leta0 = 1.69612850321655e-07 weta0 = -4.03664138925878e-22 peta0 = -1.89326617253043e-29   etab = 0.168121187844631 letab = -5.23347976377017e-08 wetab = -7.94093388050907e-23 petab = 6.31088724176809e-30   dsub = 0.859824805873 ldsub = -1.33958660221943e-7   voffl = 0.0   minv = 0.0   pclm = 1.22461387968457 lpclm = -1.36614664050484e-7   pdiblc1 = 1.20431371137557 lpdiblc1 = -2.36355661550387e-7   pdiblc2 = 0.0297230673133886 lpdiblc2 = -5.9336645927765e-9   pdiblcb = -0.075   drout = -1.12677207747957 ldrout = 4.82253601494128e-7   pscbe1 = 799984715.139714 lpscbe1 = 0.00354980180736675   pscbe2 = 7.82227156672143e-09 lpscbe2 = 3.20140480424717e-16   pvag = 0.0   delta = 0.01   alpha0 = 3.48067040171071e-08 lalpha0 = -8.06038906104501e-15   alpha1 = -3.31775714285714e-10 lalpha1 = 1.00276887212857e-16   beta0 = 38.77269915712 lbeta0 = -7.00617443553142e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.68505445252858e-11 lagidl = 1.30416208710441e-17   bgidl = 3428207740.50428 lbgidl = -563.934250277937   cgidl = -710.414937822942 lcgidl = 0.000234661796404814   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.5589   kt2 = -0.12196   at = 249570.1 lat = -0.0491356747343   ute = -0.5720187 lute = 6.31744389441e-8   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 3.7985e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.8 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.914461018033334+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.89647269488845e-8   k1 = -0.772116334006666 lk1 = 4.1671578265771e-7   k2 = 0.547754670220667 lk2 = -1.70825549075048e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 250898.039313333 lvsat = -0.0410134726498465   ua = -6.50515919813331e-10 lua = -3.71684224047192e-16   ub = 6.97168938860002e-19 lub = 3.54243188361136e-25   uc = 3.16993913027333e-13 luc = -3.76033914826469e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00776475945133333 lu0 = -8.43541285026008e-10   a0 = -1.334722697082 la0 = 4.33424125128415e-7   keta = -0.119586709834073 lketa = 2.23439889082827e-8   a1 = 0.0   a2 = -0.763969173301 la2 = 3.56649296015914e-7   ags = 1.25   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.230984759064667+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.17106883607475e-7   nfactor = {2.28364241413333+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.29495508545673e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.941101102379667 leta0 = 2.58236438351011e-7   etab = -0.324929090897333 letab = 6.21726782481684e-8   dsub = 0.438215072280667 ldsub = -3.60427508632589e-8   voffl = 0.0   minv = 0.0   pclm = 2.72696275947367 lpclm = -4.85524674939343e-7   pdiblc1 = 1.31313430735367 lpdiblc1 = -2.61628483222128e-7   pdiblc2 = 0.0294115079762267 lpdiblc2 = -5.86130711763601e-9   pdiblcb = -0.559817460262953 lpdiblcb = 1.12595461423849e-7   drout = 0.610855796801333 ldrout = 7.87016910875079e-8   pscbe1 = 894962459.092333 lpscbe1 = -22.0543663869807   pscbe2 = 1.051628577668e-08 lpscbe2 = -3.05525461738695e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 16.8847740312 lbeta0 = -1.92285704051238e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.00682062774333e-10 lagidl = -2.03622424216695e-17   bgidl = 690941011.263333 lbgidl = 71.7767867211696   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.324901909999999 lkt1 = -2.0525680698413e-7   kt2 = -0.12196   at = 38000.0   ute = -0.3   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 3.7985e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.9 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0785398795575+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.12894143648303e-8   k1 = 0.444173535962439 wk1 = -6.7238173495025e-8   k2 = 0.0137566191569487 wk2 = 2.89463132207702e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.85101710776957e-10 wua = 1.58381618737236e-16   ub = 1.08254150473868e-18 wub = -5.23004431237563e-25   uc = -7.47561310814578e-11 wuc = 5.69536897573633e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01123622823255 wu0 = -4.20882551792047e-9   a0 = 1.5598607382346 wa0 = -1.49127860082213e-6   keta = 0.0298074809386764 wketa = -1.71277283542055e-7   a1 = 0.0   a2 = 1.22113931716973 wa2 = -1.53825492252545e-6   ags = 0.0421846055410811 wags = 6.60361980738986e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.244248316605588+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 6.02621523483982e-8   nfactor = {0.78290256604464+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.7541283532912e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.556146426815906 wpclm = 3.87042084936829e-6   pdiblc1 = 0.39   pdiblc2 = 0.00986626795470871 wpdiblc2 = -4.790940083387e-8   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.01147535353239e-08 wpscbe2 = -5.12655177875429e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 0.435335040182871 wbeta0 = 2.92262781224211e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 288559453.65366 wbgidl = 6194.42081808442   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.479244701003996 wkt1 = 2.13379053251426e-7   kt2 = 0.0985606791681226 wkt2 = -7.36588456863294e-7   at = 93123.1584900001 wat = -0.0154295029170202   ute = -0.771395675491429 wute = 2.99723048747943e-6   ua1 = 7.4841500568991e-10 wua1 = 5.98247945162703e-15   ub1 = -8.77941868671241e-20 wub1 = -3.28352097100955e-24   uc1 = -6.53280162127226e-10 wuc1 = 3.78041096856005e-15   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.10 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0785398795575+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.12894143648337e-8   k1 = 0.444173535962439 wk1 = -6.72381734950266e-8   k2 = 0.0137566191569487 wk2 = 2.89463132207702e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.85101710776957e-10 wua = 1.58381618737236e-16   ub = 1.08254150473868e-18 wub = -5.23004431237566e-25   uc = -7.47561310814579e-11 wuc = 5.69536897573633e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01123622823255 wu0 = -4.2088255179205e-9   a0 = 1.5598607382346 wa0 = -1.49127860082214e-6   keta = 0.0298074809386764 wketa = -1.71277283542055e-7   a1 = 0.0   a2 = 1.22113931716973 wa2 = -1.53825492252545e-6   ags = 0.0421846055410811 wags = 6.60361980738986e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.244248316605588+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 6.02621523483991e-8   nfactor = {0.78290256604464+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.7541283532912e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.556146426815906 wpclm = 3.87042084936829e-6   pdiblc1 = 0.39   pdiblc2 = 0.00986626795470871 wpdiblc2 = -4.790940083387e-8   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.01147535353239e-08 wpscbe2 = -5.12655177875434e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 0.435335040182867 wbeta0 = 2.92262781224211e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 288559453.65366 wbgidl = 6194.42081808442   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.479244701003996 wkt1 = 2.13379053251424e-7   kt2 = 0.0985606791681226 wkt2 = -7.36588456863294e-7   at = 93123.1584899999 wat = -0.0154295029170202   ute = -0.771395675491429 wute = 2.99723048747943e-6   ua1 = 7.48415005689912e-10 wua1 = 5.98247945162703e-15   ub1 = -8.77941868671237e-20 wub1 = -3.28352097100954e-24   uc1 = -6.53280162127226e-10 wuc1 = 3.78041096856005e-15   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.11 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0807963154609+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.81693702081106e-08 wvth0 = 5.71576137410924e-08 pvth0 = 3.32702626498902e-14   k1 = 0.417796901923144 lk1 = 2.12391066806482e-07 wk1 = 1.41295662340086e-07 pk1 = -1.67916511986642e-12   k2 = 0.0215948870810933 lk2 = -6.31156380243176e-08 wk2 = -3.5911736970392e-08 pk2 = 5.22252780645434e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 276907.071027172 lvsat = -0.938847818391547 wvsat = -0.0577694330025249 pvsat = 4.6517351250855e-7   ua = -2.31585740937094e-10 lua = -2.84659649353125e-15 wua = -2.37071577384223e-15 pua = 2.03649067757163e-20   ub = 9.4342645623117e-19 lub = 1.12018817553921e-24 wub = 5.55809580010654e-25 pub = -8.68687257037535e-30   uc = -9.29749124922871e-11 luc = 1.46702055083881e-16 wuc = 1.36789595364695e-16 puc = -6.42858112075299e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0129090806374994 lu0 = -1.34702140677869e-08 wu0 = -1.64757056379129e-08 pu0 = 9.8775899578048e-14   a0 = 1.98599819919232 la0 = -3.43136238703455e-06 wa0 = -3.5309187927118e-06 pa0 = 1.64236784576623e-11   keta = 0.0728439989189316 lketa = -3.46540500650885e-07 wketa = -3.55962704849133e-07 pketa = 1.48713189092197e-12   a1 = 0.0   a2 = 1.64777902967619 la2 = -3.43540663855213e-06 wa2 = -3.09660060803028e-06 pa2 = 1.25481781376864e-11   ags = -0.129740304587892 lags = 1.38438115411165e-06 wags = 1.10524384351011e-06 pags = -3.58229686532574e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.268319362481986+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.93825910660908e-07 wvoff = 1.75943191198788e-07 pvoff = -9.31491835315764e-13   nfactor = {0.248103298835201+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.30633365579232e-06 wnfactor = 6.30646612573047e-06 pnfactor = -2.05520439617597e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.54233326552869 lpclm = 7.94101606871714e-06 wpclm = 7.67680994628947e-06 ppclm = -3.064996996096e-11   pdiblc1 = 0.39   pdiblc2 = 0.0195786608997312 lpdiblc2 = -7.82065481048066e-08 wpdiblc2 = -9.55857438701491e-08 ppdiblc2 = 3.83901499479477e-13   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.37592649480341e-08 lpscbe2 = -2.93464915114162e-14 wpscbe2 = -2.50750258693759e-14 ppscbe2 = 1.60629960856889e-19   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -3.66093372351439 lbeta0 = 3.29841514785999e-05 wbeta0 = 4.78673699090803e-05 pbeta0 = -1.50102600851485e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.50752818148432e-11 lagidl = 4.42267177533402e-16 wagidl = 2.7134745232042e-16 pagidl = -2.18495562351494e-21   bgidl = 785598093.596884 lbgidl = -4002.27590921236 wbgidl = 4017.98485304297 pbgidl = 0.0175251912644533   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.487254098726205 lkt1 = 6.44936167428696e-08 wkt1 = 3.87149318483427e-07 pkt1 = -1.39924040182252e-12   kt2 = 0.156984003677642 lkt2 = -4.70438805818505e-07 wkt2 = -1.02075623175295e-06 pkt2 = 2.28818797618084e-12   at = 93325.5382957894 lat = -0.00162961137450912 wat = -0.0380590571024162 pat = 1.82218669282477e-7   ute = -1.34458156008609 lute = 4.61543202692619e-06 wute = 6.03356519664003e-06 pute = -2.44493049074955e-11   ua1 = -4.54837732588209e-11 lua1 = 6.39266588549846e-15 wua1 = 8.79360792761429e-15 pua1 = -2.26358895928692e-20   ub1 = 3.97809371752907e-19 lub1 = -3.91019785567323e-24 wub1 = -4.82792378328722e-24 pub1 = 1.24359067343433e-29   uc1 = -1.18876329294289e-09 luc1 = 4.31184029172854e-15 wuc1 = 7.63842952118226e-15 puc1 = -3.10657028842223e-20   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.12 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08142303329579+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.07089831674929e-08 wvth0 = 4.89091365245232e-08 pvth0 = 6.66950967114026e-14   k1 = 0.515487396881226 lk1 = -1.83474557553947e-07 wk1 = -6.33612722657309e-07 pk1 = 1.46095195888057e-12   k2 = -0.0113478069284217 lk2 = 7.03761631768814e-08 wk2 = 2.29770488211215e-07 pk2 = -5.54356156571158e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 36790.0932581563 lvsat = 0.0341645239541015 wvsat = 0.11553886600505 pvsat = -2.37113828986801e-7   ua = -1.28594117381605e-09 lua = 1.42590792886446e-15 wua = 7.36450104040504e-15 pua = -1.90845574132995e-20   ub = 1.41902724578513e-18 lub = -8.07061794725304e-25 wub = -4.42252901914894e-24 pub = 1.14865651696989e-29   uc = -6.25301307791934e-11 luc = 2.33324015004685e-17 wuc = -1.29176555353035e-16 puc = 4.3490136040757e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00824054436795969 lu0 = 5.44782935070144e-09 wu0 = 2.70555253816187e-08 pu0 = -7.76232266022318e-14   a0 = 1.09551680595209 la0 = 1.77084605353388e-07 wa0 = 9.21732005951636e-07 pa0 = -1.61954457266609e-12   keta = -0.00891329850485985 lketa = -1.52400644664075e-08 wketa = 2.44006099180878e-08 pketa = -5.41926888002959e-14   a1 = 0.0   a2 = 0.8   ags = -0.0484198579680248 lags = 1.05485094353942e-06 wags = 7.03257750962221e-07 pags = -1.95335153570121e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.231301864447183+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.38220133718615e-08 wvoff = -2.74002315164229e-08 pvoff = -1.0749487402201e-13   nfactor = {0.764667236261175+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.21309105630548e-06 wnfactor = 4.98787661382106e-06 pnfactor = -1.52087988422514e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.161576664091279 leta0 = -3.30568466027235e-07 weta0 = -3.36001783376159e-14 peta0 = 1.36156087250639e-19   etab = -0.141315443783421 letab = 2.8898750786326e-07 wetab = -1.75916884683457e-16 petab = 7.12859243578084e-22   dsub = 0.86783645 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = 1.03019244767797 lpclm = -2.48348324494457e-06 wpclm = -3.92275548009014e-06 ppclm = 1.63542878411288e-11   pdiblc1 = 0.39   pdiblc2 = 0.000469570603682 lpdiblc2 = -7.71870716273331e-10 wpdiblc2 = -3.42363832267821e-09 ppdiblc2 = 1.04382524094768e-14   pdiblcb = -0.025   drout = 0.56   pscbe1 = 772293838.389157 lpscbe1 = 112.272099444406 wpscbe1 = 195.424969131564 ppscbe1 = -0.000791909463188599   pscbe2 = 5.3342763796662e-09 lpscbe2 = 4.79360943983274e-15 wpscbe2 = 2.04616743383925e-14 ppscbe2 = -2.38958138031391e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 0.91199872991433 lbeta0 = 1.44535179547205e-05 wbeta0 = 2.05251203061938e-05 pbeta0 = -3.93051612939348e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.09849436370314e-10 lagidl = -2.25437736844922e-16 wagidl = -5.4269490464084e-16 pagidl = 1.11374181918483e-21   bgidl = -851082715.158152 lbgidl = 2629.95244129958 wbgidl = 12265.9999131447 pbgidl = -0.0158977700267384   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.481199407159293 lkt1 = 3.99585352236934e-08 wkt1 = 1.02851188857615e-07 pkt1 = -2.47195296133246e-13   kt2 = 0.125626203319314 lkt2 = -3.43369378821075e-07 wkt2 = -9.08305697037346e-07 pkt2 = 1.83251108403326e-12   at = 101536.98771319 lat = -0.0349043997960257 wat = 0.0392696722591306 pat = -1.31136132971745e-7   ute = -0.326656644914016 lute = 4.90552914894544e-07 wute = 1.0501026496722e-06 pute = -4.25510368578294e-12   ua1 = 1.03635384584508e-09 lua1 = 2.00879696634803e-15 wua1 = 9.11333630151497e-15 pua1 = -2.39315066579096e-20   ub1 = -3.58794930930807e-19 lub1 = -8.44253366353275e-25 wub1 = -4.68640528085983e-24 pub1 = 1.18624393735114e-29   uc1 = 9.51813817925386e-11 luc1 = -8.91015528855392e-16 wuc1 = -2.35320271920777e-15 puc1 = 9.42281892047252e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.13 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.09992008978982+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.86694378779903e-08 wvth0 = 1.41840232409424e-07 pvth0 = -1.2402209430072e-13   k1 = 0.322318618400091 lk1 = 2.12954715902514e-07 wk1 = 2.10083151061987e-07 pk1 = -2.70516992088732e-13   k2 = 0.0714194815704112 lk2 = -9.94824252738288e-08 wk2 = -1.46926708180493e-07 pk2 = 2.18718027843351e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -77816.1399181971 lvsat = 0.269364363746641 wvsat = 0.780862922895791 pvsat = -1.60252046747243e-6   ua = -4.71190284158451e-10 lua = -2.46158881179116e-16 wua = -1.90663457852858e-15 pua = -5.79342372923273e-23   ub = 1.00523756394486e-18 lub = 4.21351833036129e-26 wub = 1.15863698142519e-24 pub = 3.26563131826077e-32   uc = -5.35895201653438e-11 luc = 4.9840959524699e-18 wuc = 7.29710923929828e-17 puc = 2.00452653543376e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0119558243997003 lu0 = -2.17682808747794e-09 wu0 = -1.24655994066535e-08 pu0 = 3.48372509662628e-15   a0 = 0.93035606372375 la0 = 5.16034582466309e-07 wa0 = 2.92354318468083e-06 pa0 = -5.72774755153484e-12   keta = -0.0731590458282234 lketa = 1.16607820757734e-07 wketa = 4.6301122191169e-07 pketa = -9.54328246989883e-13   a1 = 0.0   a2 = 0.43485314900077 la2 = 7.49370068935214e-07 wa2 = 1.80395404865712e-06 pa2 = -3.70215206867823e-12   ags = 1.50150587792378 lags = -2.12597329846438e-06 wags = -8.31569883513454e-06 pags = 1.65557389854198e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.187442773325166+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.61874993696591e-08 wvoff = -3.25029342960102e-07 pvoff = 5.03312386534494e-13   nfactor = {3.02886636110236+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.43359574825596e-06 wnfactor = -1.22289160402019e-05 pnfactor = 2.01242433644187e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.514572958182558 leta0 = 1.05705486323689e-06 weta0 = 6.72003557951116e-14 peta0 = -7.07111049841823e-20   etab = 27.1559156189137 letab = -5.57315638599394e-05 wetab = -0.000134158358467831 petab = 2.75325552057448e-10   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = -1.53054867886613 lpclm = 2.77177980681767e-06 wpclm = 1.18537845338066e-05 ppclm = -1.60230059666107e-11   pdiblc1 = 0.433359227600418 lpdiblc1 = -8.89836713283651e-08 wpdiblc1 = -1.6877794079236e-07 ppdiblc1 = 3.46373347545536e-13   pdiblc2 = -0.000260662221861173 lpdiblc2 = 7.26744488317866e-10 wpdiblc2 = 3.41211462722873e-09 ppdiblc2 = -3.59037373169904e-15   pdiblcb = -0.0505692387675422 lpdiblcb = 5.2474291276017e-08 wpdiblcb = 3.2423025342266e-10 ppdiblcb = -6.65399267975053e-16   drout = 0.646601718351473 ldrout = -1.77727770274782e-07 wdrout = -1.737288926789e-06 pdrout = 3.56533903898022e-12   pscbe1 = 855412323.221685 lpscbe1 = -58.3072292237566 wpscbe1 = -390.849938263131 ppscbe1 = 0.000411269111587811   pscbe2 = 1.85314817826693e-09 lpscbe2 = 1.1937730423257e-14 wpscbe2 = 4.92264399509419e-14 ppscbe2 = -8.29281026781344e-20   pvag = 0.0   delta = 0.01   alpha0 = -0.000163027879963663 lalpha0 = 3.34573030684568e-10 walpha0 = 8.05415639475039e-10 palpha0 = -1.65290860820317e-15   alpha1 = 4.6514685099923e-10 lalpha1 = -7.49370068935213e-16 walpha1 = -1.80395404865712e-15 palpha1 = 3.70215206867823e-21   beta0 = -69.6228909516618 lbeta0 = 0.000159208251559507 wbeta0 = 0.000381005844074919 pbeta0 = -7.79099203283235e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = -998225041.249221 lbgidl = 2931.9242500237 wbgidl = 12418.677700549 pbgidl = -0.0162111019471944   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.455768755703267 lkt1 = -1.22313412123763e-08 wkt1 = -1.70815790795682e-09 pkt1 = -3.26141086490253e-14   kt2 = -0.0366326681386286 lkt2 = -1.0374745683612e-08 wkt2 = -2.52116472603726e-08 pkt2 = 2.0187502036816e-14   at = -92117.1994361468 lat = 0.362521050201891 wat = 1.12944536540338 pat = -2.36844156799719e-6   ute = 0.304913897221569 lute = -8.05583309209416e-07 wute = -3.24755956218703e-06 pute = 4.56474350486968e-12   ua1 = 2.24395376539898e-09 lua1 = -4.6949151535703e-16 wua1 = -5.78488325572655e-15 pua1 = 6.64326014090242e-21   ub1 = -4.15783628695607e-19 lub1 = -7.27298710286347e-25 wub1 = 2.92234404183888e-24 pub1 = -3.7525631627518e-30   uc1 = -6.82764099515153e-10 luc1 = 7.05517639539947e-16 wuc1 = 4.58782675187565e-15 puc1 = -4.82186022435214e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.14 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.10111954339496+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.99315545378227e-08 wvth0 = 1.50269655689681e-07 pvth0 = -1.32891895941405e-13   k1 = 0.59576995343323 lk1 = -7.47825372267615e-08 wk1 = -2.14141723783566e-07 pk1 = 1.75870662893373e-13   k2 = -0.061070586894606 lk2 = 3.99293218380062e-08 wk2 = 1.71542997967444e-07 pk2 = -1.16389491162873e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 295848.68656071 lvsat = -0.123821834262004 wvsat = -1.53266222443628 pvsat = 8.31870174131712e-7   ua = -2.15536987707817e-10 lua = -5.15168272796219e-16 wua = -3.06468706062165e-15 pua = 1.16061838062273e-21   ub = 1.11586067652388e-18 lub = -7.42672125458617e-26 wub = 6.79331706542552e-26 pub = 1.18034176313965e-30   uc = -8.50464524643807e-11 luc = 3.80844327656054e-17 wuc = 1.70822452485754e-16 puc = -8.29181433437597e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0125253014771267 lu0 = -2.77605635586037e-09 wu0 = -1.56325665006633e-08 pu0 = 6.81614405252845e-15   a0 = 1.96395506466888 la0 = -5.71562731085193e-07 wa0 = -5.15751715019829e-06 pa0 = 2.77549161841937e-12   keta = 0.0802453961271881 lketa = -4.4810929458754e-08 wketa = -8.62960972980472e-07 pketa = 4.40916713280031e-13   a1 = 0.0   a2 = 1.53720076648239 la2 = -4.10567495126498e-07 wa2 = -3.65584555750081e-06 pa2 = 2.04288384830421e-12   ags = -1.88907118486637 lags = 1.44173768181712e-06 wags = 1.4712011186893e-05 pags = -7.67500769128851e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.13129961291441+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.05263746909754e-07 wvoff = -3.11652748066097e-07 pvoff = 4.89236958193444e-13   nfactor = {2.56258352977038+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.9429529029667e-06 wnfactor = -7.22106445700071e-07 pnfactor = 8.0162835162713e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -54.3137291937274 letab = 2.99942996066485e-05 wetab = 0.000268316125211714 petab = -1.48175406072967e-10   dsub = 0.196441259500033 ldsub = 6.68792397799072e-08 wdsub = 1.39500080652588e-07 pdsub = -1.46787983366121e-13   voffl = 0.0   minv = 0.0   pclm = 1.63638769613064 lpclm = -5.60606825218048e-07 wpclm = -7.11416470978897e-06 ppclm = 3.93588584931808e-12   pdiblc1 = 0.638319002092778 lpdiblc1 = -3.04651159319529e-07 wpdiblc1 = 7.04004558070398e-07 ppdiblc1 = -5.72005927405309e-13   pdiblc2 = 0.00043   pdiblcb = 0.247035677535084 lpdiblcb = -2.60678398669008e-07 wpdiblcb = -6.48460506845561e-10 ppdiblcb = 3.58107775681783e-16   drout = -0.0991772767029468 ldrout = 6.07012956818266e-07 wdrout = 3.47457785357799e-06 pdrout = -1.91881129759347e-12   pscbe1 = 800000000.0   pscbe2 = -4.55099964314322e-09 lpscbe2 = 1.8676450139301e-14 wpscbe2 = 9.19873252036396e-14 ppscbe2 = -1.27922944859089e-19   pvag = 0.0   delta = 0.01   alpha0 = 0.000326056059927326 lalpha0 = -1.80062121478147e-10 walpha0 = -1.61083127895008e-09 palpha0 = 8.89570297981229e-16   alpha1 = -6.3029370199846e-10 lalpha1 = 4.03299584872736e-16 walpha1 = 3.60790809731424e-15 palpha1 = -1.99244199138511e-21   beta0 = 161.535400990813 lbeta0 = -8.40264430289184e-05 wbeta0 = -0.000756558405281379 pbeta0 = 4.17894815152184e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 3194920884.18433 lbgidl = -1480.28419799228 wbgidl = -10133.9143846545 pbgidl = 0.00751970520631641   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.422034696479698 lkt1 = -4.7727768891962e-08 wkt1 = -6.88230117011279e-08 pkt1 = 3.80070264508664e-14   kt2 = -0.036888055239614 lkt2 = -1.01060163943099e-08 wkt2 = -1.26825546227599e-08 pkt2 = 7.00385201253676e-15   at = 437105.801160867 lat = -0.194350147615313 wat = -2.28196819870442 pat = 1.2211944749403e-6   ute = -0.41698182272101 lute = -4.59735911698759e-08 wute = 1.29867374002565e-06 pute = -2.18998663750498e-13   ua1 = 3.25359550859553e-09 lua1 = -1.5318799721434e-15 wua1 = 1.30166634692508e-15 pua1 = -8.13512072640545e-22   ub1 = -2.69245915495752e-18 lub1 = 1.66831717549407e-24 wub1 = -2.00248830881652e-24 pub1 = 1.4295572043989e-30   uc1 = -5.26933091723513e-11 luc1 = 4.25300608972668e-17 wuc1 = 1.12967210435006e-17 puc1 = -6.23853511922593e-24   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.15 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.98905946004674+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.95284207065057e-09 wvth0 = -2.33244481469658e-07 pvth0 = 7.89011017058809e-14   k1 = 0.0161666531471547 lk1 = 2.45299328133122e-07 wk1 = 2.57139904214025e-07 pk1 = -8.43913171969013e-14   k2 = 0.171374220713287 lk2 = -8.84366960497995e-08 wk2 = -1.41438253747832e-07 pk2 = 5.64522142281266e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 34737.0375707444 lvsat = 0.0203752461111616 wvsat = 0.221597406356101 pvsat = -1.36907427155965e-7   ua = -2.01904558056641e-10 lua = -5.22696686644072e-16 wua = -1.55436727117142e-15 pua = 3.26554849137364e-22   ub = -2.01063387760547e-19 lub = 6.5299488348676e-25 wub = 4.569910975776e-24 pub = -1.3058439658942e-30   uc = -3.55763345787711e-11 luc = 1.07649064541027e-17 wuc = 4.52001529218703e-17 puc = -1.3544107765702e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0101610037596452 lu0 = -1.47038949146522e-09 wu0 = -2.89175711221637e-09 pu0 = -2.19878746575658e-16   a0 = 1.29956995977867 la0 = -2.04660707605311e-07 wa0 = -5.67591168252314e-07 pa0 = 2.40737124371582e-13   keta = 0.0400587508168046 lketa = -2.26181358926118e-08 wketa = 2.53191981866346e-07 pketa = -1.75470942963441e-13   a1 = 0.0   a2 = 0.786185871032144 la2 = 4.17522378163174e-09 wa2 = 9.58749203731416e-08 pa2 = -2.89775235583396e-14   ags = -0.241731280691576 lags = 5.32005751115915e-07 wags = -2.64878007239631e-06 pags = 1.91236775611517e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.420940952436176+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.46886553517641e-08 wvoff = 1.12798219043705e-06 pvoff = -3.05791359150348e-13   nfactor = {-6.0772198847667+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.8283180540875e-06 wnfactor = 3.78490645332388e-05 pnfactor = -1.32843756586508e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 2.33326720822035 leta0 = -1.01793141286923e-06 weta0 = -8.69556302967029e-06 peta0 = 4.80206381419421e-12   etab = 0.0165841055287816 letab = -9.2356006726557e-09 wetab = -7.38230302812677e-08 petab = 4.10641140372919e-14   dsub = 0.211319899988026 ldsub = 5.86626147208963e-08 wdsub = -3.72966792547118e-07 pdsub = 1.36218260090305e-13   voffl = 0.0   minv = 0.0   pclm = 0.196965973173891 lpclm = 2.34303745332755e-07 wpclm = 1.70309381075847e-06 ppclm = -9.33383447844613e-13   pdiblc1 = -0.481128527581577 lpdiblc1 = 3.13555902810426e-07 wpdiblc1 = 3.91396554750628e-07 ppdiblc1 = -3.99370345827991e-13   pdiblc2 = -0.0216592707351792 lpdiblc2 = 1.21986451386076e-08 wpdiblc2 = 7.22451168577391e-08 ppdiblc2 = -3.98968600688685e-14   pdiblcb = -0.25702711300154 lpdiblcb = 1.76867489653095e-08 wpdiblcb = -1.03632427781087e-06 ppdiblcb = 5.7230282815111e-13   drout = 2.47632903292781 ldrout = -8.15292374131156e-07 wdrout = -5.78919447767648e-06 pdrout = 3.1970421259355e-12   pscbe1 = 800014851.523919 lpscbe1 = -0.00820165012373764 wpscbe1 = -0.0733717588700529 ppscbe1 = 4.0519040234166e-8   pscbe2 = 6.8382533994105e-08 lpscbe2 = -2.16005832771339e-14 wpscbe2 = -4.08902049159795e-13 ppscbe2 = 1.48689705907498e-19   pvag = 0.0   delta = 0.01   alpha0 = -8.50482994908932e-09 lalpha0 = 4.75195710557493e-15 walpha0 = -7.72493941457803e-15 palpha0 = 4.26604371712481e-21   alpha1 = 2.208972e-10 lalpha1 = -6.67646324196e-17   beta0 = 1.93829072440572 lbeta0 = 4.10994393593332e-06 wbeta0 = -1.04123648005583e-07 pbeta0 = 1.48233300125103e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = -147626182.901117 lbgidl = 365.614021976192 wbgidl = 3495.13804975464 pbgidl = -6.84359721903234e-6   cgidl = 502.446090441154 lcgidl = -0.000111799436323494 wcgidl = 0.000558490781082388 pcgidl = -3.08422624417282e-10   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.47465545335372 lkt1 = -1.8668324253582e-08 wkt1 = 1.88611018561579e-07 pkt1 = -1.04159114723502e-13   kt2 = 0.0364676062722873 lkt2 = -5.06161669746267e-08 wkt2 = -7.58589371357557e-08 pkt2 = 4.18925670206612e-14   at = 2341.23036150483 lat = 0.0457455432566399 wat = 0.403589153950563 pat = -2.61885774161948e-7   ute = -0.47799715396112 lute = -1.22783015998442e-08 wute = 6.86970683808241e-07 pute = 1.18810067124172e-13   ua1 = 9.97351018687055e-10 lua1 = -2.85884746302872e-16 wua1 = -1.07635728068468e-15 pua1 = 4.9973482954155e-22   ub1 = 2.97854444586369e-19 lub1 = 1.69374223411532e-26 wub1 = 9.69175125004363e-25 pub1 = -2.1152312528465e-31   uc1 = -6.05646700353748e-11 luc1 = 4.68769648343455e-17 wuc1 = 4.7447070735293e-16 puc1 = -2.62023126840704e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.16 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.981508510571743+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.23506369282269e-09 wvth0 = 3.66179920463012e-08 pvth0 = -2.66294187700318e-15   k1 = 0.288093281588083 lk1 = 1.63111408173249e-07 wk1 = -8.26846886346771e-07 pk1 = 2.43236102342565e-13   k2 = 0.0689686861092151 lk2 = -5.74853400544609e-08 wk2 = 4.08487525666276e-07 pk2 = -1.09759003119332e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 194867.00986066 lvsat = -0.0280229171036593 wvsat = -1.00122351950783 pvsat = 2.32681637939926e-7   ua = -7.62797261216702e-10 lua = -3.53170793362865e-16 wua = -2.79617897790234e-15 pua = 7.01883744814845e-22   ub = 3.52545968344313e-19 lub = 4.85670330869559e-25 wub = 6.17214820846123e-24 pub = -1.79010895381268e-30   uc = 1.87015446872389e-13 luc = -4.43157476978569e-20 wuc = -1.98242315929724e-18 puc = 7.16495576798345e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00697988579148386 lu0 = -5.08918853414227e-10 wu0 = -5.2273957769716e-10 pu0 = -9.3589771326133e-16   a0 = 0.824195115181821 la0 = -6.09819884498251e-08 wa0 = 1.68117047134461e-06 pa0 = -4.38935339865112e-13   keta = -0.283869466253851 lketa = 7.52869002194742e-08 wketa = 5.28306336081656e-08 pketa = -1.14913127981844e-13   a1 = 0.0   a2 = 0.808410646650161 la2 = -2.5420590754848e-09 wa2 = 5.93187087269924e-07 pa2 = -1.79286644817725e-13   ags = 2.4091487663693 lags = -2.69204186947906e-07 wags = 1.58827502956271e-05 pags = -3.68865757690731e-12   b0 = 0.0   b1 = 1.72706074707307e-23 lb1 = -5.21992021377607e-30 wb1 = -1.19864098554822e-28 pb1 = 3.62280847395052e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.0832924883662316+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -9.77123724966781e-08 wvoff = -9.75991759290343e-07 pvoff = 3.30120039337107e-13   nfactor = {8.56199269541531+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.59628147378445e-06 wnfactor = -3.08380880765288e-05 pnfactor = 7.47583540758314e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -4.81391124640607 leta0 = 1.14225324479242e-06 weta0 = 2.95270946192026e-05 peta0 = -6.75046690157407e-12   etab = 0.141427327376964 letab = -4.6968590573716e-08 wetab = 1.85264793223264e-07 petab = -3.72433670021884e-14   dsub = 0.976112258175267 ldsub = -1.7249052199469e-07 wdsub = -8.07075875418434e-07 pdsub = 2.67424691624581e-13   voffl = 0.0   minv = 0.0   pclm = 2.0972640620747 lpclm = -3.40048049950891e-07 wpclm = -6.05649961318172e-06 ppclm = 1.41189934738734e-12   pdiblc1 = 1.81689140471563 lpdiblc1 = -3.81004535586879e-07 wpdiblc1 = -4.2515049416436e-06 ppdiblc1 = 1.00391413114669e-12   pdiblc2 = 0.0672676998180687 lpdiblc2 = -1.46789092223177e-08 wpdiblc2 = -2.60572972802049e-07 ppdiblc2 = 6.06950778041748e-14   pdiblcb = -0.608281024994499 lpdiblcb = 1.23850785087798e-07 wpdiblcb = 3.70115813503883e-06 ppdiblcb = -8.59568068755823e-13   drout = -4.42034835135399 ldrout = 1.26918008852633e-06 wdrout = 2.28585793382521e-05 pdrout = -5.46154697551222e-12   pscbe1 = 799946958.843145 lpscbe1 = 0.0123184373919685 wpscbe1 = 0.262041995956679 ppscbe1 = -6.0857419267174e-8   pscbe2 = -4.25072845052935e-08 lpscbe2 = 1.19150881355799e-14 wpscbe2 = 3.49304845209432e-13 ppscbe2 = -8.04730204673408e-20   pvag = 0.0   delta = 0.01   alpha0 = 3.08315355324619e-08 lalpha0 = -7.13718400666553e-15 walpha0 = 2.75890693377786e-14 palpha0 = -6.40736823021371e-21   alpha1 = -3.31775714285714e-10 lalpha1 = 1.00276887212857e-16   beta0 = 38.3514677573478 lbeta0 = -6.89568393003418e-06 wbeta0 = 2.9234942721184e-06 pbeta0 = -7.66843022906862e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -4.97362091163676e-11 lagidl = 4.52567210519583e-17 wagidl = 7.39749610127707e-16 pagidl = -2.23584141413828e-22   bgidl = 2031246879.15712 lbgidl = -292.935108919475 wbgidl = 9695.40038736469 pbgidl = -0.0018808294869253   cgidl = -423.02175157555 lcgidl = 0.00016791674065116 wcgidl = -0.0019946099324371 pcgidl = 4.6323419453899e-10   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.53642139749 wkt1 = -1.56009418383204e-7   kt2 = -0.131000844526 wkt2 = 6.27466451958831e-8   at = 662440.426151353 lat = -0.153764817976471 wat = -2.86546547641926 pat = 7.26163104484919e-7   ute = -1.24395279149307 lute = 2.19226428154725e-07 wute = 4.66345925014893e-06 pute = -1.08305576663234e-12   ua1 = -2.24384786026297e-10 lua1 = 8.33763485211055e-17 wua1 = 2.49161965650814e-15 pua1 = -5.7866122388642e-22   ub1 = 2.25143101946728e-19 lub1 = 3.8913916674586e-26 wub1 = 1.1629038860292e-24 pub1 = -2.7007628720308e-31   uc1 = 9.45322712812e-11 wuc1 = -3.92457978640474e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.17 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.730495956357789+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.25309723211339e-08 wvth0 = -1.27678232052301e-06 pvth0 = 3.02365086915034e-13   k1 = -0.956662217122414 lk1 = 4.52197159460272e-07 wk1 = 1.28081342588331e-06 pk1 = -2.46253251550685e-13   k2 = 0.612962051445456 lk2 = -1.83823991200246e-07 wk2 = -4.52562191739707e-07 pk2 = 9.02137664001849e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 399779.037998857 lvsat = -0.0756123012545586 wvsat = -1.03328656676527 pvsat = 2.40128056224137e-7   ua = -1.01584061719131e-09 lua = -2.94403245241257e-16 wua = 2.53548206716152e-15 pua = -5.36357211273917e-22   ub = 1.89532010524645e-18 lub = 1.27371836992999e-25 wub = -8.31559108356268e-24 pub = 1.57456708258483e-30   uc = -7.75201567193427e-13 luc = 1.7915241829983e-19 wuc = 7.58022130398021e-18 puc = -1.5043616612866e-24   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00899922352002942 lu0 = -9.77895905504839e-10 wu0 = -8.56761541499581e-09 pu0 = 9.3246838582042e-16   a0 = 1.3614730004898 la0 = -1.85761016367407e-07 wa0 = -1.8712547741273e-05 pa0 = 4.29736295898784e-12   keta = 0.361083192452804 lketa = -7.44988400965354e-08 wketa = -3.33601841381052e-06 pketa = 6.72123341337814e-13   a1 = 0.0   a2 = -3.36873416813813 la2 = 9.67570584145393e-07 wa2 = 1.80779864624009e-05 pa2 = -4.24000890609627e-12   ags = 1.25   b0 = 0.0   b1 = -4.02980840983717e-23 lb1 = 8.15000542230699e-30 wb1 = 2.79682896627919e-28 pb1 = -5.65639080627203e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.654648500672143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.3040580686264e-07 wvoff = -2.94037558112568e-06 pvoff = 7.8633443127161e-13   nfactor = {0.0694583730429557+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.76050174846272e-07 wnfactor = 1.53672170807865e-05 pnfactor = -3.25502327806721e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -2.15914687284473 leta0 = 5.25702802383416e-07 weta0 = 8.45366664274789e-06 peta0 = -1.8563107680383e-12   etab = -0.301609313190094 letab = 5.59235679414993e-08 wetab = -1.6184747051395e-07 petab = 4.33710264649339e-14   dsub = 0.054051239356947 ldsub = 4.16516951987327e-08 wdsub = 2.66623230299256e-06 pdsub = -5.39226819654125e-13   voffl = 0.0   minv = 0.0   pclm = 4.93771199806277 lpclm = -9.99722199948568e-07 wpclm = -1.53433783416902e-05 ppclm = 3.56871192393233e-12   pdiblc1 = 1.23373547982464 lpdiblc1 = -2.45570654122421e-07 wpdiblc1 = 5.51055827318498e-07 ppdiblc1 = -1.11446989519373e-13   pdiblc2 = 0.0459169913146829 lpdiblc2 = -9.72035662736592e-09 wpdiblc2 = -1.14553867600118e-07 ppdiblc2 = 2.67831627547629e-14   pdiblcb = -1.7574019634672 lpdiblcb = 3.90726079201513e-07 wpdiblcb = 8.3116582414995e-06 ppdiblcb = -1.93032444498057e-12   drout = 1.34473754542752 ldrout = -6.97207553998973e-08 wdrout = -5.0933978086176e-06 pdrout = 1.03010405300825e-12   pscbe1 = 1129536455.93944 lpscbe1 = -76.5325351367437 wpscbe1 = -1628.02615508063 ppscbe1 = 0.00037809767833439   pscbe2 = 1.25199286412875e-08 lpscbe2 = -8.64596927221575e-16 wpscbe2 = -1.39059871633932e-14 ppscbe2 = 3.88015287542127e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 22.6573581293564 lbeta0 = -3.25083682770058e-06 wbeta0 = -4.00637667453247e-05 pbeta0 = 9.21664743756712e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1023242628185e-09 lagidl = -2.22301259131611e-16 wagidl = -6.25771442668938e-15 pagidl = 1.40152789888868e-21   bgidl = -1853663781.65044 lbgidl = 609.308197678453 wbgidl = 17660.4534726296 pbgidl = -0.00373065731060649   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.448960930258432 lkt1 = -2.28848147943279e-07 wkt1 = -8.61013294180471e-07 pkt1 = 1.63732215126783e-13   kt2 = -0.19194909517506 lkt2 = 1.41548045754897e-08 wkt2 = 4.85748970674241e-07 pkt2 = -9.82393290760704e-14   at = -253430.002860088 lat = 0.0589396780684328 wat = 2.02262686149602 pat = -4.09062124349539e-7   ute = -0.3   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 4.75741930805324e-10 luc1 = -8.85332749568611e-17 wuc1 = -3.03818727777998e-15 puc1 = 6.14452109620056e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.18 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0779365737308+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.8308871096619e-8   k1 = 0.44163999375501 wk1 = -5.47215826767618e-8   k2 = 0.0188717449284315 wk2 = 3.6757903623484e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 317436.83559945 wvsat = -0.776249557052281   ua = -1.08568402148447e-09 wua = 2.63143453872216e-15   ub = 1.42006531196265e-18 wub = -2.1904909148089e-24   uc = -1.12127974134718e-11 wuc = -2.56972758524605e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00931695215140001 wu0 = 5.27307429199628e-9   a0 = 1.3885541675039 wa0 = -6.4496380723826e-7   keta = -0.0120162226354518 wketa = 3.53465424225372e-8   a1 = 0.0   a2 = 1.07116081478027 wa2 = -7.97308298292954e-7   ags = 0.233117095552106 wags = -2.82911766338459e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.237524997059419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 2.70465858371805e-8   nfactor = {1.28514856689764+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.27285621803587e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.342711317998797 wpclm = -5.70252987714072e-7   pdiblc1 = 0.39   pdiblc2 = 0.000134606789153327 wpdiblc2 = 1.68432815036079e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 863028978.109892 wpscbe1 = -311.385350668957   pscbe2 = 7.90654360323031e-09 wpscbe2 = 5.78278301732606e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.20825201062161e-10 walpha0 = -5.96919047882889e-16   alpha1 = 2.47017517295807e-10 walpha1 = -7.26318315010878e-16   beta0 = 1.45762335603557 wbeta0 = 2.41758137921639e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1821530357.50449 wbgidl = -1378.99535929101   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.423900194041174 wkt1 = -6.00423034802669e-8   kt2 = -0.0474057316515528 wkt2 = -1.54629780442067e-8   at = 90000.0   ute = -0.155112624558572 wute = -4.74248390194267e-8   ua1 = 1.73808613484057e-09 wua1 = 1.09315551145107e-15   ub1 = -7.7294082115852e-19 wub1 = 1.01344711034548e-25   uc1 = 1.1389025772369e-10 wuc1 = -9.68110292534689e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.19 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0779365737308+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.8308871096619e-8   k1 = 0.44163999375501 wk1 = -5.47215826767618e-8   k2 = 0.0188717449284315 wk2 = 3.6757903623484e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 317436.83559945 wvsat = -0.776249557052281   ua = -1.08568402148447e-09 wua = 2.63143453872216e-15   ub = 1.42006531196265e-18 wub = -2.1904909148089e-24   uc = -1.12127974134718e-11 wuc = -2.56972758524605e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0093169521514 wu0 = 5.27307429199624e-9   a0 = 1.3885541675039 wa0 = -6.44963807238262e-7   keta = -0.0120162226354518 wketa = 3.53465424225372e-8   a1 = 0.0   a2 = 1.07116081478027 wa2 = -7.97308298292952e-7   ags = 0.233117095552106 wags = -2.82911766338459e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.237524997059419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 2.70465858371805e-8   nfactor = {1.28514856689764+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.27285621803587e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.342711317998797 wpclm = -5.70252987714072e-7   pdiblc1 = 0.39   pdiblc2 = 0.000134606789153327 wpdiblc2 = 1.68432815036079e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 863028978.109891 wpscbe1 = -311.385350668957   pscbe2 = 7.9065436032303e-09 wpscbe2 = 5.78278301732606e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.20825201062161e-10 walpha0 = -5.96919047882889e-16   alpha1 = 2.47017517295807e-10 walpha1 = -7.26318315010878e-16   beta0 = 1.45762335603557 wbeta0 = 2.41758137921639e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1821530357.50449 wbgidl = -1378.99535929101   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.423900194041174 wkt1 = -6.00423034802669e-8   kt2 = -0.0474057316515528 wkt2 = -1.54629780442067e-8   at = 90000.0   ute = -0.155112624558572 wute = -4.74248390194269e-8   ua1 = 1.73808613484057e-09 wua1 = 1.09315551145107e-15   ub1 = -7.7294082115852e-19 wub1 = 1.01344711034549e-25   uc1 = 1.1389025772369e-10 wuc1 = -9.68110292534689e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.20 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.079655991715+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.38451714273555e-08 wvth0 = 5.15240128143245e-08 pvth0 = 5.46333276095941e-14   k1 = 0.52902793972395 lk1 = -7.03668976212774e-07 wk1 = -4.08224839967412e-07 pk1 = 2.84649412899584e-12   k2 = -0.0138018187073352 lk2 = 2.63095474071157e-07 wk2 = 1.38960456344224e-07 pk2 = -1.08934500465989e-12   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 541388.299083055 lvsat = -1.80331160417562 wvsat = -1.36439984988711 pvsat = 4.7359290784272e-6   ua = -1.61701905226823e-09 lua = 4.27843878228337e-15 wua = 4.47381273374584e-15 pua = -1.4835276924232e-20   ub = 1.81495069936404e-18 lub = -3.17971309650513e-24 wub = -3.74982713190414e-24 pub = 1.25561541387517e-29   uc = 3.61721922968067e-12 luc = -1.19414897704708e-16 wuc = -3.40409555090618e-16 puc = 6.71853361091102e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00742805119970565 lu0 = 1.52098894659742e-08 wu0 = 1.06025102033561e-08 pu0 = -4.29139130111961e-14   a0 = 1.38691933667273 la0 = 1.31640551164983e-08 wa0 = -5.7125821628963e-07 pa0 = -5.93495328776973e-13   keta = -0.0124902349173079 lketa = 3.81686207849022e-09 wketa = 6.56184650190479e-08 pketa = -2.43756876824295e-13   a1 = 0.0   a2 = 1.34586319317218 la2 = -2.2119703034896e-06 wa2 = -1.60503004094284e-06 pa2 = 6.50397174820032e-12   ags = 0.278648108189909 lags = -3.66626777795659e-07 wags = -9.12338750011207e-07 pags = 5.06829902329e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.240658345913799+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.52304863792353e-08 wvoff = 3.92880271419035e-08 pvoff = -9.85710600558706e-14   nfactor = {1.18324602555231+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.20544025230134e-07 wnfactor = 1.68653169847959e-06 pnfactor = -3.33101549167452e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.202964430553487 lpclm = 1.12527589620329e-06 wpclm = -9.45575366205042e-07 ppclm = 3.02218699494726e-12   pdiblc1 = 0.39   pdiblc2 = 0.000322175716321631 lpdiblc2 = -1.51035058080849e-09 wpdiblc2 = -4.51924930024346e-10 ppdiblc2 = 4.99527131015859e-15   pdiblcb = -0.025   drout = 0.56   pscbe1 = 926881161.945632 lpscbe1 = -514.153300326056 wpscbe1 = -626.837627556664 ppscbe1 = 0.0025400983884031   pscbe2 = 6.39572520032322e-09 lpscbe2 = 1.21654769090798e-14 wpscbe2 = 1.13034539230152e-14 ppscbe2 = -4.44537836556388e-20   pvag = 0.0   delta = 0.01   alpha0 = 2.15976674931938e-10 lalpha0 = 3.90415105924054e-17 walpha0 = -5.72965621148684e-16 palpha0 = -1.92878812746514e-22   alpha1 = 2.483361246689e-10 lalpha1 = -1.0617746989733e-17 walpha1 = -7.32832699847472e-16 palpha1 = 5.24554096997708e-23   beta0 = -9.28893859359682 lbeta0 = 8.65339282329937e-05 wbeta0 = 7.56716961506028e-05 pbeta0 = -4.14657358249563e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.53228408002491e-10 lagidl = -4.28608075739201e-16 wagidl = -2.62967082577604e-16 pagidl = 2.11747484991593e-21   bgidl = 1436019384.2205 lbgidl = 3104.2280360492 wbgidl = 804.674598983758 pbgidl = -0.0175834411358283   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.369529976334523 lkt1 = -4.37802204936857e-07 wkt1 = -1.94449308567387e-07 pkt1 = 1.08227786586372e-12   kt2 = -0.0433313336730128 lkt2 = -3.28080426019123e-08 wkt2 = -3.11279141789043e-08 pkt2 = 1.26137872336066e-13   at = 14131.695244995 lat = 0.610910025885356 wat = 0.353186419640031 pat = -2.8439428752415e-6   ute = -0.0295059265910812 lute = -1.01141565446184e-06 wute = -4.63371602463442e-07 pute = 3.34930441431473e-12   ua1 = 1.28904040780381e-09 lua1 = 3.61582531221167e-15 wua1 = 2.20058845374833e-15 pua1 = -8.91731915758251e-21   ub1 = -6.20728708040466e-19 lub1 = -1.22564892237006e-24 wub1 = 2.04013060003741e-25 pub1 = -8.26710494308739e-31   uc1 = 3.61312057858612e-10 luc1 = -1.99230045818383e-15 wuc1 = -1.94886483157261e-17 puc1 = 7.89727387168625e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.21 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08582799843499+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.88556424543794e-08 wvth0 = 7.06712157409009e-08 pvth0 = -2.29557914192004e-14   k1 = 0.374091023629722 lk1 = -7.58269425283502e-08 wk1 = 6.49351610077834e-08 pk1 = 9.29134827164106e-13   k2 = 0.0443847484234683 lk2 = 2.73093647213288e-08 wk2 = -4.55679642331161e-08 pk2 = -3.41591004074312e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 96946.613403905 lvsat = -0.00232589447407894 wvsat = -0.181655530641344 pvsat = -5.68383100262196e-8   ua = 1.5316884201651e-10 lua = -2.89479272101673e-15 wua = 2.54790707644622e-16 pua = 2.26122554788244e-21   ub = 5.18699296725806e-19 lub = 2.07301257607583e-24 wub = 2.54081447078062e-26 pub = -2.74201658425216e-30   uc = -6.24672366597151e-11 luc = 1.48375376081905e-16 wuc = -1.29487274454567e-16 puc = -1.82854974160372e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0140174043478232 lu0 = -1.14917707030132e-08 wu0 = -1.48419752899208e-09 pu0 = 6.06436379025764e-15   a0 = 1.30089108880114 la0 = 3.61771420356412e-07 wa0 = -9.28892841450629e-08 pa0 = -2.53196248547725e-12   keta = -0.0138206242705174 lketa = 9.207923022308e-09 wketa = 4.8644527560571e-08 pketa = -1.74974357575744e-13   a1 = 0.0   a2 = 0.8   ags = 0.107430152800773 lags = 3.27189983404277e-07 wags = -6.66961926094333e-08 pags = 1.64154988955656e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.228238471803584+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.50978615447635e-08 wvoff = -4.25344701026908e-08 pvoff = 2.32993581646057e-13   nfactor = {1.8045916860669+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.69729957817049e-06 wnfactor = -1.49716429610439e-07 pnfactor = 4.1099081316414e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.281508709155915 leta0 = -8.16562256116094e-07 weta0 = -5.92506576285756e-07 peta0 = 2.40098062620792e-12   etab = -0.246161704882658 letab = 7.13850035478817e-07 wetab = 5.17977456507474e-07 petab = -2.09897052229022e-12   dsub = 1.32041024149884 ldsub = -3.081367078242e-06 wdsub = -2.23587392649366e-06 pdsub = 9.06030446751645e-12   voffl = 0.0   minv = 0.0   pclm = -0.0187617362594414 lpclm = 2.02376420358781e-06 wpclm = 1.25944763022428e-06 ppclm = -5.91310200717249e-12   pdiblc1 = 0.39   pdiblc2 = -0.000867984940361258 lpdiblc2 = 3.31246960911015e-09 wpdiblc2 = 3.18435715195809e-09 ppdiblc2 = -9.73982730258018e-15   pdiblcb = 0.0106965096431757 lpdiblcb = -1.44650931325991e-07 wpdiblcb = -1.76353329947984e-07 ppdiblcb = 7.1462654680841e-13   drout = 0.56   pscbe1 = 829273386.331941 lpscbe1 = -118.622874849902 wpscbe1 = -86.0740659025705 ppscbe1 = 0.000348793031035237   pscbe2 = 8.70320199564189e-09 lpscbe2 = 2.81502021758724e-15 wpscbe2 = 3.81799525987074e-15 ppscbe2 = -1.41208861861224e-20   pvag = 0.0   delta = 0.01   alpha0 = 2.79727693131376e-10 lalpha0 = -2.19293106649142e-16 walpha0 = -8.8791810416252e-16 palpha0 = 1.08338518187892e-21   alpha1 = 3.95238137923471e-10 lalpha1 = -6.05900401886478e-16 walpha1 = -1.45858038421412e-15 palpha1 = 2.99336138344075e-21   beta0 = 13.4101560631088 lbeta0 = -5.44831919597901e-06 wbeta0 = -4.12201787707996e-05 pbeta0 = 5.90169236575655e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 8.24178752175675e-11 lagidl = -1.41666589935225e-16 wagidl = 8.68618888495646e-17 pagidl = 6.99882849252988e-22   bgidl = 2560499674.46556 lbgidl = -1452.43934873431 wbgidl = -4588.41865091409 pbgidl = 0.00427068323441749   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.504256596664946 lkt1 = 1.08142799210759e-07 wkt1 = 2.16761825757691e-07 pkt1 = -5.84049574727132e-13   kt2 = -0.075427424620915 lkt2 = 9.72531172690874e-08 wkt2 = 8.49700360751479e-08 pkt2 = -3.44319233895266e-13   at = 173540.552996234 lat = -0.0350534020750983 wat = -0.316453299894799 pat = -1.30400009234522e-7   ute = -1.39801352356609 lute = 4.53410967582696e-06 wute = 6.34298296210611e-06 pute = -2.42316982254803e-11   ua1 = 3.53644749639054e-10 lua1 = 7.4062758202402e-15 wua1 = 1.24861596869164e-14 pua1 = -5.05969531881893e-20   ub1 = 4.4777817981316e-19 lub1 = -5.5554984791267e-24 wub1 = -8.67116052298463e-24 pub1 = 3.51376495311408e-29   uc1 = -5.37989394832776e-10 luc1 = 1.65188755837468e-15 wuc1 = 7.74883920068803e-16 puc1 = -3.14001794091137e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.22 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0773601454227+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.1477550384889e-08 wvth0 = 3.03861616234483e-08 pvth0 = 5.97189288979653e-14   k1 = 0.0965716161820174 lk1 = 4.93710318770349e-07 wk1 = 1.32535285011345e-06 pk1 = -1.65754855237917e-12   k2 = 0.147995848085386 lk2 = -1.85325789282145e-07 wk2 = -5.25240928960757e-07 pk2 = 6.42814480077236e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 232573.684212345 lvsat = -0.280665601151204 wvsat = -0.752572127605146 pvsat = 1.11482127967656e-6   ua = -1.78728053355777e-09 lua = 1.08748092685996e-15 wua = 4.5953147804899e-15 pua = -6.64658459694576e-21   ub = 1.8781255819182e-18 lub = -7.16860501726265e-25 wub = -3.15373725852302e-24 pub = 3.78236231551048e-30   uc = 5.21831304723287e-11 luc = -8.69150373122623e-17 wuc = -4.49583054884674e-16 puc = 4.7405935055685e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0064415963943534 lu0 = 4.05562813883955e-09 wu0 = 1.47766290508636e-08 pu0 = -2.7306803732465e-14   a0 = 2.47321129186457 la0 = -2.0441145101391e-06 wa0 = -4.69870503594617e-06 pa0 = 6.9202906504463e-12   keta = 0.10428461487845 lketa = -2.33172727284487e-07 wketa = -4.13622957636578e-07 pketa = 7.73710853047709e-13   a1 = 0.0   a2 = 0.8   ags = -1.15266060776887 lags = 2.913202426148e-06 wags = 4.79681840162339e-06 pags = -8.33956389185559e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.314431375247064+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.51790921196794e-07 wvoff = 3.02339075919668e-07 pvoff = -4.74770739063507e-13   nfactor = {-1.31780174744975+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.71061048901001e-06 wnfactor = 9.24515531255331e-06 pnfactor = -1.5170651637112e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.754437048311831 leta0 = 1.30945017302679e-06 weta0 = 1.18501315257151e-06 peta0 = -1.24692179470131e-12   etab = -35.0184112517041 letab = 7.20749557621962e-05 wetab = 0.000173004714070945 petab = -3.56083668332113e-10   dsub = -0.64514758299769 ldsub = 9.52435208176239e-07 wdsub = 4.47174785298732e-06 pdsub = -4.70536537607094e-12   voffl = 0.0   minv = 0.0   pclm = 1.86165589263554 lpclm = -1.83530971238852e-06 wpclm = -4.9049007838617e-06 ppclm = 6.73763887519657e-12   pdiblc1 = 0.391214694947652 lpdiblc1 = -2.49284920345284e-09 wpdiblc1 = 3.94308938167068e-08 ppdiblc1 = -8.09217758190803e-14   pdiblc2 = 0.00107868910114834 lpdiblc2 = -6.82578565859638e-10 wpdiblc2 = -3.20475262797425e-09 ppdiblc2 = 3.37217851951751e-15   pdiblcb = -0.121919018695504 lpdiblcb = 1.27508358398365e-07 wpdiblcb = 3.52817272490044e-07 ppdiblcb = -3.71360117850817e-13   drout = 0.213762113279117 ldrout = 7.10564279357725e-07 wdrout = 4.01091168377354e-07 pdrout = -8.23136542664244e-13   pscbe1 = 741453227.336118 lpscbe1 = 61.6054317081607 wpscbe1 = 172.148131805145 ppscbe1 = -0.000181141666655041   pscbe2 = 1.33333377790773e-08 lpscbe2 = -6.68714353301769e-15 wpscbe2 = -7.48973999983892e-15 ppscbe2 = 9.08533434646995e-21   pvag = 0.0   delta = 0.01   alpha0 = 2.49551793485874e-10 lalpha0 = -1.57364827832956e-16 walpha0 = -7.38838531961881e-16 palpha0 = 7.77437673387165e-22   alpha1 = 1.0e-10   beta0 = 12.5926840823319 lbeta0 = -3.77066804573347e-06 wbeta0 = -2.51680529185366e-05 pbeta0 = 2.60740607421395e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -7.77493824450987e-11 lagidl = 1.87035543432178e-16 wagidl = 8.78144552611285e-16 pagidl = -9.24021458473356e-22   bgidl = 2580327557.44461 lbgidl = -1493.13098278289 wbgidl = -5260.63250322379 pbgidl = 0.00565022940732311   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.39015704202572 lkt1 = -1.26017213100712e-07 wkt1 = -3.25853131920598e-07 pkt1 = 5.29528173863433e-13   kt2 = -0.0111784209943443 lkt2 = -3.46014506805168e-08 wkt2 = -1.50964593138981e-07 pkt2 = 1.39875957367026e-13   at = 355265.45570987 lat = -0.407997061594839 wat = -1.08078251918908 pat = 1.43818928075763e-6   ute = 1.65928818671363 lute = -1.74021635798263e-06 wute = -9.93864556290258e-06 pute = 9.18215994356911e-12   ua1 = 3.5712495972144e-09 lua1 = 8.02968795037629e-16 wua1 = -1.23421921384867e-14 pua1 = 3.5685804703147e-22   ub1 = -6.27644511410636e-19 lub1 = -3.3484697890215e-24 wub1 = 3.96901141985401e-24 pub1 = 9.1969451426538e-30   uc1 = 7.23011429834593e-10 luc1 = -9.35992557043153e-16 wuc1 = -2.35719947725353e-15 puc1 = 3.28777828665961e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.23 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.09620926030654+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.13113995775971e-08 wvth0 = 1.26011127831141e-07 pvth0 = -4.09017724193146e-14   k1 = 0.608889241138781 lk1 = -4.53723158670304e-08 wk1 = -2.78955625662116e-07 pk1 = 3.05738110963376e-14   k2 = -0.0444713314397418 lk2 = 1.71964531029145e-08 wk2 = 8.95368297626435e-08 pk2 = -4.0811130951512e-15   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -166376.105993038 lvsat = 0.139126522943878 wvsat = 0.750891046351173 pvsat = -4.67187320876756e-7   ua = 1.3774111491287e-10 lua = -9.38109627591731e-16 wua = -4.81000531211559e-15 pua = 3.25009763325772e-21   ub = 6.28569889043862e-19 lub = 5.97975729210909e-25 wub = 2.47532128462088e-24 pub = -2.14077513310289e-30   uc = -4.31700842475558e-11 luc = 1.34197154042332e-17 wuc = -3.60615553622471e-17 puc = 3.89342473348738e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0140900582680962 lu0 = -3.99241232857319e-09 wu0 = -2.33630161553942e-08 pu0 = 1.28253709583034e-14   a0 = 0.286902736168719 la0 = 2.56413363431969e-07 wa0 = 3.12771201042259e-06 pa0 = -1.3150019016759e-12   keta = -0.228911781264145 lketa = 1.17430848181786e-07 wketa = 6.64384368490593e-07 pketa = -3.60614809818324e-13   a1 = 0.0   a2 = 0.859980227324859 la2 = -6.31137743409914e-08 wa2 = -3.10137576988722e-07 pa2 = 3.26340094423344e-13   ags = 2.61023367141765 lags = -1.04627673886606e-06 wags = -7.51613945832053e-06 pags = 4.61665982556538e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.139871384391731+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.18886072607941e-08 wvoff = -2.6930517799022e-07 pvoff = 1.26737925603396e-13   nfactor = {4.33176556322851+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.23410716668e-06 wnfactor = -9.46248879689542e-06 pnfactor = 4.51433592354671e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 70.453484032735 letab = -3.89071077475878e-05 wetab = -0.000348077851139509 petab = 1.92221813332631e-10   dsub = 0.220369307733666 ldsub = 4.17011185224044e-08 wdsub = 2.12870949198516e-08 pdsub = -2.23991966197498e-14   voffl = 0.0   minv = 0.0   pclm = -0.443483944051648 lpclm = 5.90257544786719e-07 wpclm = 3.16113372350319e-06 ppclm = -1.74978947293659e-12   pdiblc1 = 1.07222161960949 lpdiblc1 = -7.190776186304e-07 wpdiblc1 = -1.43962719296405e-06 ppdiblc1 = 1.47540674258936e-12   pdiblc2 = 0.000685606979147342 lpdiblc2 = -2.68960654558937e-10 wpdiblc2 = -1.26278850176592e-09 ppdiblc2 = 1.32876036146368e-15   pdiblcb = 0.246949198818305 lpdiblcb = -2.60630641403017e-07 wpdiblcb = -2.21225188150361e-10 ppdiblcb = 1.2217006157947e-16   drout = 0.766501933441765 ldrout = 1.28947672770319e-07 wdrout = -8.02182336754706e-07 pdrout = 4.42999580196429e-13   pscbe1 = 800000000.0   pscbe2 = 2.70962484782613e-08 lpscbe2 = -2.11690699758591e-14 wpscbe2 = -6.43612266768871e-14 ppscbe2 = 6.89279581019871e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.51748137307525 lbeta0 = 5.17435478662877e-07 wbeta0 = -5.9598945846429e-07 pbeta0 = 2.18278970722649e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.74653096206734e-10 lagidl = -1.83777497911863e-16 wagidl = -8.62847808081751e-16 pagidl = 9.07925566119367e-22   bgidl = 740971024.204828 lbgidl = 442.31905382294 wbgidl = 1989.46220478488 pbgidl = -0.00197863199851605   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.511527507385962 lkt1 = 1.69400948134563e-09 wkt1 = 3.73302993543815e-07 pkt1 = -2.06153965063618e-13   kt2 = -0.0317733584777374 lkt2 = -1.29305718781789e-08 wkt2 = -3.795095802263e-08 pkt2 = 2.09581509112913e-14   at = -141757.546284682 lat = 0.114991913092915 wat = 0.577820613347566 pat = -3.07064255232127e-7   ute = 0.362333931118972 lute = -3.75505321212935e-07 wute = -2.55142055895237e-06 pute = 1.40900414373753e-12   ua1 = 8.81074951395768e-09 lua1 = -4.71025831585607e-15 wua1 = -2.61526316692046e-14 pua1 = 1.48887963701527e-20   ub1 = -8.56010681760827e-18 lub1 = 4.99840814543881e-24 wub1 = 2.69857577301849e-23 pub1 = -1.50222650451677e-29   uc1 = -3.77278781679422e-10 luc1 = 2.21780115990989e-16 wuc1 = 1.61486327423185e-15 puc1 = -8.91796939151619e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.24 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.04869165024445+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.50701320440791e-08 wvth0 = 6.1359540564396e-08 pvth0 = -5.19838591236848e-15   k1 = 0.0748214304123809 lk1 = 2.49562894131949e-07 wk1 = -3.26353536887455e-08 pk1 = -1.0545483485905e-13   k2 = 0.134378963210011 lk2 = -8.15723701653488e-08 wk2 = 4.13313480480453e-08 pk2 = 2.25400267433637e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160099.697218241 lvsat = -0.0411674540489278 wvsat = -0.397738285031259 pvsat = 1.67135186973873e-7   ua = -7.47475709297361e-10 lua = -4.49254832939399e-16 wua = 1.1409463661172e-15 pua = -3.62737743845909e-23   ub = 1.07647164937017e-18 lub = 3.50625117383028e-25 wub = -1.74156205548981e-24 pub = 1.87969173289862e-31   uc = -5.34728965500016e-11 luc = 1.91093713785727e-17 wuc = 1.33615472228875e-16 puc = -5.47687034131303e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00971904382758901 lu0 = -1.57855020090418e-09 wu0 = -7.08319389570716e-10 pu0 = 3.14473252254692e-16   a0 = 0.552548889412001 la0 = 1.0971213482644e-07 wa0 = 3.12295602018001e-06 pa0 = -1.31237543935637e-12   keta = 0.128797135047934 lketa = -8.01113968891451e-08 wketa = -1.85206889894358e-07 pketa = 1.08566015485956e-13   a1 = 0.0   a2 = 0.680039545350283 la2 = 3.62572076946946e-08 wa2 = 6.20275153977444e-07 pa2 = -1.87473823363605e-13   ags = -3.5696135284376 lags = 2.3665006183236e-06 wags = 1.37921303115967e-05 pags = -7.15068299698303e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.186289866777605+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -6.25432529257144e-09 wvoff = -3.12768168286602e-08 pvoff = -4.71157064954776e-15   nfactor = {2.18566332275233+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -4.89372270927214e-08 wnfactor = -2.97248869937096e-06 pnfactor = 9.30278799689506e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.34506864980239 leta0 = 8.00373236271787e-08 weta0 = 1.1268380924467e-06 peta0 = -6.22288448687044e-13   etab = 0.0054783332518165 letab = -2.68973608813714e-09 wetab = -1.89566037800642e-08 petab = 8.72523753626354e-15   dsub = 0.287939864256969 ldsub = 4.38575167630572e-09 wdsub = -7.51496401587114e-07 pdsub = 4.04365079841747e-13   voffl = 0.0   minv = 0.0   pclm = 0.824497345591899 lpclm = -1.09976246549903e-07 wpclm = -1.39713218553585e-06 ppclm = 7.6748096746886e-13   pdiblc1 = -0.918791677213391 lpdiblc1 = 3.80445537446958e-07 wpdiblc1 = 2.55360665889309e-06 ppdiblc1 = -7.29828699461779e-13   pdiblc2 = -0.00547892670232925 lpdiblc2 = 3.13535991930074e-09 wpdiblc2 = -7.69148138170804e-09 ppdiblc2 = 4.87896100356155e-15   pdiblcb = -0.644099910401411 lpdiblcb = 2.31444991819806e-07 wpdiblcb = 8.75951668383731e-07 ppdiblcb = -4.83738177203237e-13   drout = 1.01619461569169 ldrout = -8.94336315342509e-09 wdrout = 1.42438380281173e-06 pdrout = -7.86605984416159e-13   pscbe1 = 800000000.0   pscbe2 = -4.94128792732774e-08 lpscbe2 = 2.10825602610339e-14 wpscbe2 = 1.73048779925628e-13 ppscbe2 = -6.21800561742054e-20   pvag = 0.0   delta = 0.01   alpha0 = -2.50179149920936e-08 lalpha0 = 1.38711927289788e-14 walpha0 = 7.38555166064155e-14 palpha0 = -4.07861920572767e-20   alpha1 = 3.9863737399692e-10 lalpha1 = -1.64920399328181e-16 walpha1 = -8.78099059634066e-16 palpha1 = 4.84924058989495e-22   beta0 = -9.8874350487505 lbeta0 = 1.06814217382012e-05 wbeta0 = 5.83191266920034e-05 pbeta0 = -3.23171815175601e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.12823984538031e-09 lagidl = -2.31189380503573e-15 wagidl = -1.99009235822523e-14 pagidl = 1.14215696458746e-20   bgidl = -87269743.8592463 lbgidl = 899.709220300949 wbgidl = 3196.95598334997 pbgidl = -0.00264546198527218   cgidl = 654.130172571928 lcgidl = -0.000195565908891639 wcgidl = -0.000190882007777359 pcgidl = 1.05413252620992e-10   egidl = 2.34998158035639 legidl = -1.24253657788075e-06 wegidl = -1.11157014504731e-05 pegidl = 6.13856831611364e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.376383854291642 lkt1 = -7.29381269344209e-08 wkt1 = -2.96885292062277e-07 pkt1 = 1.63952824344348e-13   kt2 = 0.123217261218271 lkt2 = -9.85230566709614e-08 wkt2 = -5.04432785797386e-07 pkt2 = 2.78569474927106e-13   at = 67552.7518438692 lat = -0.000598233876490745 wat = 0.0814212703298167 pat = -3.29311928459767e-8   ute = -0.33894417636 lute = 1.17706046955756e-8   ua1 = 4.7802947231179e-10 lua1 = -1.08572001897423e-16 wua1 = 1.48927406345777e-15 pua1 = -3.7625257736995e-22   ub1 = 5.62917068794566e-19 lub1 = -3.97179346599469e-26 wub1 = -3.40327593640372e-25 pub1 = 6.83742923175191e-32   uc1 = 9.71610105740937e-12 luc1 = 8.06490096375307e-18 wuc1 = 1.27258945266997e-16 puc1 = -7.02778617110821e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.25 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.967256330198797+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -9.54312339247856e-09 wvth0 = -3.37927986139802e-08 pvth0 = 2.35607425379221e-14   k1 = 0.466954512139257 lk1 = 1.31043415111573e-07 wk1 = -1.71048436019494e-06 pk1 = 4.01663282414401e-13   k2 = 0.0326968128005891 lk2 = -5.0839651979154e-08 wk2 = 5.87683354764668e-07 pk2 = -1.42591042822689e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -97969.7185813092 lvsat = 0.0368322203905757 wvsat = 0.445493056091258 pvsat = -8.77255832610198e-8   ua = -2.09368685405575e-09 lua = -4.23719379141922e-17 wua = 3.77888435003708e-15 pua = -8.33572064458489e-22   ub = 2.37530890121131e-18 lub = -4.19393501251933e-26 wub = -3.82101309700666e-24 pub = 8.16468694431039e-31   uc = 4.15408143492957e-11 luc = -9.60785764476359e-18 wuc = -2.06284754545242e-16 puc = 4.79637608277592e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00585193961963768 lu0 = -4.09745023780349e-10 wu0 = 5.04971177386462e-09 pu0 = -1.4258513606755e-15   a0 = 4.04221810030529 la0 = -9.45015956481581e-07 wa0 = -1.42169964628607e-05 pa0 = 3.9285038189753e-12   keta = -0.0689173248107162 lketa = -2.03535853980871e-08 wketa = -1.00910865126513e-06 pketa = 3.57584555547944e-13   a1 = 0.0   a2 = 0.492424568336084 la2 = 9.29625211923977e-08 wa2 = 2.15426960443826e-06 pa2 = -6.51112908054233e-13   ags = 14.2472309521148 lags = -3.018515908012e-06 wags = -4.26015450745015e-05 pags = 9.89391063273744e-12   b0 = 0.0   b1 = -1.72706074707307e-23 lb1 = 5.21992021377607e-30 wb1 = 5.07816686718996e-29 pb1 = -1.53484038844009e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0890122418054879+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.56558064970192e-08 wvoff = -1.24745706516081e-07 pvoff = 2.35387469762473e-14   nfactor = {1.7275670266576+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 8.95191717278401e-08 wnfactor = 2.92638181185484e-06 pnfactor = -8.52613520234911e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.90091531339766 leta0 = -3.90206439517848e-07 weta0 = -3.64651354814226e-06 peta0 = 8.20423671219485e-13   etab = 0.0601141213568998 letab = -1.92030205923819e-08 wetab = 5.86980669473545e-07 petab = -1.74415061743727e-13   dsub = 0.147079752519742 ldsub = 4.69597344281004e-08 wdsub = 3.28863668776835e-06 pdsub = -8.16736865484316e-13   voffl = 0.0   minv = 0.0   pclm = -0.160142800373233 lpclm = 1.87624345087037e-07 wpclm = 5.09588534600802e-06 ppclm = -1.19498813031755e-12   pdiblc1 = 0.7863668039552 lpdiblc1 = -1.3492667737688e-07 wpdiblc1 = 8.39649536877311e-07 ppdiblc1 = -2.11797157032364e-13   pdiblc2 = 0.00620205011479454 lpdiblc2 = -3.95133556837204e-10 wpdiblc2 = 4.11128440539515e-08 ppdiblc2 = -9.87180472908849e-15   pdiblcb = 1.13900481561019 lpdiblcb = -3.07485929884119e-07 wpdiblcb = -4.93104931162142e-06 ppdiblcb = 1.27138721999646e-12   drout = 1.66864914059586 ldrout = -2.06143176124037e-07 wdrout = -7.22321281689679e-06 pdrout = 1.8270695607144e-12   pscbe1 = 800000000.0   pscbe2 = 5.73089260768228e-08 lpscbe2 = -1.11733583533965e-14 wpscbe2 = -1.43822390335589e-13 ppscbe2 = 3.35920369390555e-20   pvag = 0.0   delta = 0.01   alpha0 = 8.98068392574773e-08 lalpha0 = -2.08337854696743e-14 walpha0 = -2.6376970216577e-13 palpha0 = 6.12586669400849e-20   alpha1 = -9.66562049988999e-10 lalpha1 = 2.47701570175595e-16 walpha1 = 3.13606807012167e-15 palpha1 = -7.28329856809266e-22   beta0 = 81.4108197610566 lbeta0 = -1.69128366902793e-05 wbeta0 = -0.000209804870129979 pbeta0 = 4.87214196539064e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.45508960108606e-08 lagidl = 3.3337442535621e-15 wagidl = 7.23805863392265e-14 pagidl = -1.64698707573229e-20   bgidl = 8395061587.77585 lbgidl = -1664.01604836644 wbgidl = -21744.0856087522 pbgidl = 0.00489279324864956   cgidl = -964.750616328312 lcgidl = 0.000293729477387936 wcgidl = 0.000681721456347714 pcgidl = -1.58325036186562e-10   egidl = -7.93564850127281 legidl = 1.8662231148811e-06 wegidl = 3.96989337516898e-05 pegidl = -9.2197994712937e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.928951877812266 lkt1 = 9.40716901985232e-08 wkt1 = 1.78322940364396e-06 pkt1 = -4.64747281629992e-13   kt2 = -0.50081169376885 lkt2 = 9.00853267712108e-08 wkt2 = 1.88974248783666e-06 pkt2 = -4.4505324230187e-13   at = 180033.67904651 lat = -0.0345948067569986 wat = -0.482206242065008 pat = 1.37421277382772e-7   ute = -0.3   ua1 = 6.63501034644162e-11 lua1 = 1.58552055811136e-17 wua1 = 1.05528690559594e-15 pua1 = -2.45082996816318e-22   ub1 = 5.60256898053273e-19 lub1 = -3.89139166745862e-26 wub1 = -4.92676293816114e-25 pub1 = 1.14420620504736e-31   uc1 = 3.6399600638055e-11 wuc1 = -1.05262111336736e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.26 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.18409126572727+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 4.08152725394613e-08 wvth0 = 9.64138264030202e-07 pvth0 = -2.08201761243749e-13   k1 = -0.481175103572284 lk1 = 3.51239881453269e-07 wk1 = -1.06826038161571e-06 pk1 = 2.52511258957227e-13   k2 = 0.461779772627692 lk2 = -1.5049116581828e-07 wk2 = 2.94331512018645e-07 pk2 = -7.44621308078242e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -13227.6274067492 lvsat = 0.0171514629099223 wvsat = 1.00711182128598 pvsat = -2.18157610146138e-7   ua = -4.23610973820067e-10 lua = -4.30235370567767e-16 wua = -3.90340954372784e-16 pua = 1.34701327913569e-22   ub = 1.78073375870087e-19 lub = 4.68353219986627e-25 wub = 1.68212573854546e-25 pub = -1.10001043046779e-31   uc = 9.55774579715881e-13 luc = -1.82266253557053e-19 wuc = -9.71410511550707e-19 puc = 2.81173869342632e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00834687136243835 lu0 = -9.89175456523607e-10 wu0 = -5.34476599806606e-09 pu0 = 9.88193340511003e-16   a0 = -7.7099802569944 la0 = 1.78434984661277e-06 wa0 = 2.61036263165362e-05 pa0 = -5.43567857718018e-12   keta = -0.906843864304083 lketa = 1.74248987913471e-07 wketa = 2.9279878104779e-06 pketa = -5.56778538016643e-13   a1 = 0.0   a2 = 2.97695343317024 la2 = -4.84051915963282e-07 wa2 = -1.32719452392356e-05 pa2 = 2.93151750588513e-12   ags = 1.25   b0 = 0.0   b1 = 4.02980840983718e-23 lb1 = -8.150005422307e-30 wb1 = -1.18490560234432e-28 pb1 = 2.39638863734923e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0907522151314133+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.52517098718865e-08 wvoff = 7.42166485075997e-07 pvoff = -1.77795541135671e-13   nfactor = {4.92060080979784+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -6.52040573169998e-07 wnfactor = -8.59913512914887e-06 pnfactor = 1.82410711069462e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.100052773978913 leta0 = 2.80312792243812e-08 weta0 = -2.70757530267651e-06 peta0 = 6.02361836277783e-13   etab = -0.0718703584633695 letab = 1.1449450954517e-08 wetab = -1.29683882092382e-06 petab = 2.63088828164629e-13   dsub = 0.951159913084759 ldsub = -1.39782254302001e-07 wdsub = -1.76580050689772e-06 pdsub = 3.57120791916515e-13   voffl = 0.0   minv = 0.0   pclm = 1.73948772884229 lpclm = -2.53551547909564e-07 wpclm = 4.5697596284658e-07 ppclm = -1.17633898443993e-13   pdiblc1 = 1.45859139326137 lpdiblc1 = -2.91046132671113e-07 wpdiblc1 = -5.59811579311653e-07 ppdiblc1 = 1.13217890974709e-13   pdiblc2 = 0.0145784545020842 lpdiblc2 = -2.34049484095452e-09 wpdiblc2 = 4.02695416867848e-08 ppdiblc2 = -9.6759536574306e-15   pdiblcb = -0.183543633855276 lpdiblcb = -3.33310334910044e-10 wpdiblcb = 5.36243780312909e-07 ppdiblcb = 1.64667044635568e-15   drout = -0.695136458821075 ldrout = 3.42829482841351e-07 wdrout = 4.98429821599476e-06 pdrout = -1.00803942409743e-12   pscbe1 = 800000000.0   pscbe2 = 1.08502851150172e-08 lpscbe2 = -3.83664200503821e-16 wpscbe2 = -5.65736009516754e-15 ppscbe2 = 1.5041758209293e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 11.4438481180933 lbeta0 = -6.63497295002605e-07 wbeta0 = 1.5334922108541e-05 pbeta0 = -3.56572111494425e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.14643221956541e-09 lagidl = 2.20651369280327e-16 wagidl = 4.85193460832023e-15 pagidl = -7.86814093382021e-22   bgidl = 2781174665.44629 lbgidl = -360.230107863854 wbgidl = -5237.28084612927 pbgidl = 0.00105920339016372   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.596295086326148 lkt1 = -2.60156240493875e-07 wkt1 = -1.58889591624474e-06 pkt1 = 3.18405219036919e-13   kt2 = -0.0519709048249393 lkt2 = -1.41548045754898e-08 wkt2 = -2.05792589973999e-07 pkt2 = 4.16201107741115e-14   at = -15615.9678066636 lat = 0.0108434541771231 wat = 0.847741770228957 pat = -1.71449838836415e-7   ute = -0.3   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 2.57117365327937e-11 luc1 = 2.48218162339821e-18 wuc1 = -8.14879617439256e-16 puc1 = 1.64803698469768e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.27 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.058106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020121864   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.9074547e-10   ub = 6.7508962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111103   a0 = 1.169205   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.13690013   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22832658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.718041+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.28 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.058106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020121864   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.9074547e-10   ub = 6.7508962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111103   a0 = 1.169205   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.13690013   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22832658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.718041+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.29 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06213291648125+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.24257100477313e-8   k1 = 0.390192585249268 lk1 = 2.64410333808601e-7   k2 = 0.0334579811031172 lk2 = -1.07385655590756e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 77362.3059087988 lvsat = -0.192644324783984   ua = -9.54963130039224e-11 lua = -7.66969357677566e-16   ub = 5.3965206952502e-19 lub = 1.09057606774931e-24   uc = -1.12154474749911e-10 luc = 1.09079281016842e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01103391521945 lu0 = 6.15068814490277e-10   a0 = 1.1926370951475 la0 = -1.88680924126792e-7   keta = 0.00982629744199512 lketa = -7.90837090926421e-08 wketa = -3.05022850878929e-24 pketa = 1.33120277756046e-29   a1 = 0.0   a2 = 0.8   ags = -0.0316340240020127 lags = 1.35707796182363e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.227296672049727+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -8.29306908322664e-9   nfactor = {1.75682755040487+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.12318728991801e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.118621319005712 lpclm = 2.15310752635537e-06 ppclm = -8.07793566946316e-28   pdiblc1 = 0.39   pdiblc2 = 0.0001684781660675 lpdiblc2 = 1.88517775900135e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 713696623.18301 lpscbe1 = 349.722254583012   pscbe2 = 1.02399768933739e-08 lpscbe2 = -2.95304653026833e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.1113753017793e-11 lalpha0 = -2.65556694823196e-17   alpha1 = -8.96841316424275e-13 lalpha1 = 7.22209195873409e-18 walpha1 = 1.72562570700712e-34 palpha1 = 1.36067201924711e-39   beta0 = 16.4466505479362 lbeta0 = -5.44890955563207e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37945359045825e-11 lagidl = 2.91535194824077e-16   bgidl = 1709685443.33537 lbgidl = -2875.81786995767   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.435661274676058 lkt1 = -6.97245760515383e-8   kt2 = -0.0539177913697828 lkt2 = 1.00908564946196e-8   at = 134248.740964903 lat = -0.35630161469345   ute = -0.18709643648423 lute = 1.27667076618715e-7   ua1 = 2.03745022542645e-09 lua1 = 5.83086867619045e-16   ub1 = -5.5134482266655e-19 lub1 = -1.50680928618931e-24   uc1 = 3.54684059921588e-10 luc1 = -1.9654421999395e-15 wuc1 = 1.97215226305253e-31 puc1 = -7.52316384526264e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.30 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0617930492405+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.10484854004685e-8   k1 = 0.396175167497855 lk1 = 2.4016745676984e-7   k2 = 0.0288872973925624 lk2 = -8.88641345194464e-08 pk2 = 5.04870979341448e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 35166.4189627955 lvsat = -0.0216563372782503   ua = 2.39821967327356e-10 lua = -2.12576051192203e-15 pua = 7.52316384526264e-37   ub = 5.27340487637496e-19 lub = 1.14046558927195e-24   uc = -1.06505251716063e-10 luc = 8.61872565224955e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01351263572555 lu0 = -9.4293090053099e-9   a0 = 1.269299878692 la0 = -4.99337152105506e-7   keta = 0.0027231515263313 lketa = -5.03000357779147e-8   a1 = 0.0   a2 = 0.8   ags = 0.0847470903399452 lags = 8.85473405899229e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.242704245700565+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.41421633903642e-8   nfactor = {1.7536738301684+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.99539088239589e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.409570498982405 lpclm = 1.27459292557421e-8   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -0.0492804311967633 lpdiblcb = 9.83902073540655e-8   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.00016842862568e-08 lpscbe2 = -1.98742698112673e-15 wpscbe2 = 1.26217744835362e-29   pvag = 0.0   delta = 0.01   alpha0 = -2.2249091881834e-11 lalpha0 = 1.4916111522228e-16 palpha0 = 9.4039548065783e-38   alpha1 = -1.00818213493928e-10 lalpha1 = 4.1212777291542e-16 walpha1 = 3.08148791101958e-33 palpha1 = 9.99170198198944e-38   beta0 = -0.608633512779299 lbeta0 = 1.46230598917253e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.11959196440775e-10 lagidl = 9.63602863189145e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.430536915819335 lkt1 = -9.04897233581801e-8   kt2 = -0.0465295136580215 lkt2 = -1.98482401449211e-8   at = 65916.269111195 lat = -0.0794018339515661   ute = 0.759205248425275 lute = -3.70697730194403e-06 wute = 2.11758236813575e-22 pute = 1.61558713389263e-27   ua1 = 4.6001291289309e-09 lua1 = -9.80151078035453e-15 pua1 = -6.01853107621011e-36   ub1 = -2.50124286704804e-18 lub1 = 6.39465141486927e-24 pub1 = 2.80259692864963e-45   uc1 = -2.74455005969835e-10 luc1 = 5.83982175845552e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.31 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.067025954293+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.17876781641302e-8   k1 = 0.5473179077703 lk1 = -7.00141739551044e-8   k2 = -0.0306361297303179 lk2 = 3.32924021294949e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -23372.568622654 lvsat = 0.0984798902210754   ua = -2.24435517749833e-10 lua = -1.17299133797476e-15   ub = 8.0555432378014e-19 lub = 5.69503191545063e-25   uc = -1.00717959024594e-10 luc = 7.43103256074759e-17 puc = -9.4039548065783e-38   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0114670586675 lu0 = -5.2312878069662e-9   a0 = 0.875203734829 la0 = 3.09443900464329e-7   keta = -0.0363866141112533 lketa = 2.99627069834588e-8   a1 = 0.0   a2 = 0.8   ags = 0.47871484501648 lags = 7.69558391385944e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21160727277401+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.67638161934739e-9   nfactor = {1.8264322366809+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.48857018696022e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.35141963 leta0 = 8.8537791573009e-07 weta0 = 2.11758236813575e-22   etab = 23.819681025454 letab = -4.90274306567208e-05 wetab = 1.05879118406788e-21 petab = -1.4641258400902e-26   dsub = 0.8756729 ldsub = -6.478374993147e-07 pdsub = 8.07793566946316e-28   voffl = 0.0   minv = 0.0   pclm = 0.19352212829884 lpclm = 4.56129685652493e-7   pdiblc1 = 0.40462495709812 lpdiblc1 = -3.00139658299168e-8   pdiblc2 = -1.12322449999998e-05 lpdiblc2 = 4.64283541175535e-10   pdiblcb = -0.00192751819088942 lpdiblcb = 1.21052310815198e-9   drout = 0.35017133948588 ldrout = 4.3061939973948e-7   pscbe1 = 800000000.0   pscbe2 = 1.07861123141011e-08 lpscbe2 = -3.59726391027389e-15   pvag = 0.0   delta = 0.01   alpha0 = -1.72372784857094e-12 lalpha0 = 1.07038080562564e-16   alpha1 = 1.0e-10   beta0 = 4.0331472627167 lbeta0 = 5.09699778767909e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.2090346350012e-10 lagidl = -1.27219823143757e-16   bgidl = 791211102.8839 lbgidl = 428.485552584237   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.50097816472 lkt1 = 5.40728366094671e-8   kt2 = -0.062520771458 lkt2 = 1.29697067362804e-8   at = -12303.612781 lat = 0.0811243711225178   ute = -1.72079858075 lute = 1.38259319645412e-06 pute = 1.61558713389263e-27   ua1 = -6.2627209372e-10 lua1 = 9.24334544022214e-16 pua1 = -3.76158192263132e-37   ub1 = 7.2219766731e-19 lub1 = -2.20631857683276e-25   uc1 = -7.8661062751e-11 luc1 = 1.82165426432301e-16 wuc1 = 2.46519032881566e-32 puc1 = 9.4039548065783e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.32 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.053353466422+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.74008985092845e-8   k1 = 0.51401774048586 lk1 = -3.49743060312228e-8   k2 = -0.014020275351072 lk2 = 1.58084856699141e-08 wk2 = -4.96308367531817e-24 pk2 = 1.57772181044202e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 88998.418987736 lvsat = -0.0197616948950443 wvsat = 1.11022302462516e-16   ua = -1.4981191443158e-09 lua = 1.6723334229389e-16   ub = 1.4704150546063e-18 lub = -1.30091858441647e-25   uc = -5.54344501838022e-11 luc = 2.66610704143146e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00614440599032001 lu0 = 3.69436214027714e-10   a0 = 1.350622929424 la0 = -1.90812619113898e-07 wa0 = -1.6940658945086e-21   keta = -0.0029577719143154 lketa = -5.21255821637372e-9   a1 = 0.0   a2 = 0.75450389119454 la2 = 4.78729620177834e-8   ags = 0.0540298743621399 lags = 5.23827626714829e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.23146081302896+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.12143671391419e-8   nfactor = {1.1136174798474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.01197319478732e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -47.9261614871143 letab = 2.64666299062316e-5   dsub = 0.22760894893034 ldsub = 3.40832567506922e-8   voffl = 0.0   minv = 0.0   pclm = 0.63160281715444 lpclm = -4.83765263098929e-9   pdiblc1 = 0.5826111596911 lpdiblc1 = -2.17298701604962e-7   pdiblc2 = 0.00025613852915488 lpdiblc2 = 1.82944515666482e-10   pdiblcb = 0.246873961168832 lpdiblcb = -2.60589091937759e-07 wpdiblcb = -3.63959469523332e-23 ppdiblcb = -8.83524213847533e-29   drout = 0.49368348102824 ldrout = 2.79609753386521e-7   pscbe1 = 800000000.0   pscbe2 = 5.207296985686e-09 lpscbe2 = 2.27300546734361e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.3147881520168 lbeta0 = 5.91671133399287e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.879739862914e-11 lagidl = 1.25003731125722e-16   bgidl = 1417577794.2322 lbgidl = -230.604413820173   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.38456890918 lkt1 = -6.84179876677095e-8   kt2 = -0.044680301402 lkt2 = -5.8028029968553e-9   at = 54756.535718 lat = 0.0105607992854845   ute = -0.50539224092 lute = 1.03690383212383e-7   ua1 = -8.36379234399999e-11 lua1 = 3.53351536784276e-16 pua1 = 1.88079096131566e-37   ub1 = 6.1762288776e-19 lub1 = -1.10593777925246e-25 wub1 = -7.3468396926393e-40   uc1 = 1.7192864804e-10 luc1 = -8.15158426195538e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.33 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.027823558128+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.33021853632811e-8   k1 = 0.0637222996046001 lk1 = 2.13698199127367e-7   k2 = 0.148435560935972 lk2 = -7.3906612728752e-08 wk2 = -2.64697796016969e-23 pk2 = 1.89326617253043e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24830.77092048 lvsat = 0.0156744395765614   ua = -3.594451984908e-10 lua = -4.61591373570345e-16   ub = 4.841745580592e-19 lub = 4.14552552093013e-25   uc = -8.030900781986e-12 luc = 4.82792082007395e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00947814772352 lu0 = -1.47159932193985e-9   a0 = 1.61465159268 la0 = -3.36620600196381e-7   keta = 0.065809139972256 lketa = -4.31886039373496e-08 wketa = -2.64697796016969e-23 pketa = -6.31088724176809e-30   a1 = 0.0   a2 = 0.89099221761092 la2 = -2.75017608273773e-8   ags = 1.121025338429 lags = -6.54131493478461e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.19692696556756+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -7.85670838448397e-9   nfactor = {1.1747338499596+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.67446231898861e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.72830100286768 leta0 = -1.31600060726656e-07 weta0 = 8.470329472543e-22   etab = -0.000968718832646104 letab = 2.77676297448353e-10   dsub = 0.0323594607981201 ldsub = 1.41908419825294e-7   voffl = 0.0   minv = 0.0   pclm = 0.34933923849988 lpclm = 1.51040432835941e-7   pdiblc1 = -0.0503220228321601 lpdiblc1 = 1.3223421791123e-7   pdiblc2 = -0.00809476346559456 lpdiblc2 = 4.7946716859529e-09 ppdiblc2 = 1.18329135783152e-30   pdiblcb = -0.3461928541026 lpdiblcb = 6.69279053281821e-8   drout = 1.50062087007432 ldrout = -2.76464371152453e-7   pscbe1 = 800000000.0   pscbe2 = 9.44019959449479e-09 lpscbe2 = -6.45853680527897e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.94662656196521 lbeta0 = -3.09500205625848e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.63997097720492e-09 lagidl = 1.57252849167915e-15 wagidl = -1.18329135783152e-30 pagidl = 1.88079096131566e-37   bgidl = 1000000000.0   cgidl = 589.212096506972 lcgidl = -0.0001597153558113   egidl = -1.4304163768928 legidl = 8.45161731224411e-07 pegidl = 3.53409685539013e-28   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.47735315044 lkt1 = -1.71785399215632e-8   kt2 = -0.048337964648 lkt2 = -3.78288407289453e-9   at = 95243.744212 lat = -0.0117979781948675 wat = 1.11022302462516e-16   ute = -0.33894417636 lute = 1.17706046955755e-8   ua1 = 9.8452460016e-10 lua1 = -2.36533739736159e-16   ub1 = 4.4717324952e-19 lub1 = -1.64641583546734e-26   uc1 = 5.29962718026e-11 luc1 = -1.58362703690832e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.34 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.978749102599998+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.53022529886812e-9   k1 = -0.114773200682 lk1 = 2.67647214620489e-7   k2 = 0.232565166926557 lk2 = -9.93341972321643e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53540.3814982856 lvsat = 0.00699716074669365   ua = -8.0850600053857e-10 lua = -3.25865889577021e-16   ub = 1.07580025833286e-18 lub = 2.35737825565202e-25   uc = -2.86156636893698e-11 luc = 6.70439257742381e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00756932292285713 lu0 = -8.9467038771311e-10   a0 = -0.792915753 la0 = 3.91049777063979e-7   keta = -0.412110446799685 lketa = 1.01259245727362e-07 pketa = -5.04870979341448e-29   a1 = 0.0   a2 = 1.225081562433 la2 = -1.28477926674437e-7   ags = -0.241354828357858 lags = 3.46356719402314e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.131437671832571+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.76503889908281e-8   nfactor = {2.72281576313714+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -2.0045068978566e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.660753149102428 leta0 = -1.11184194761085e-7   etab = 0.25974349550927 letab = -7.85207655018953e-08 wetab = -7.83753630393994e-23 petab = -1.16356983520099e-29   dsub = 1.26552967418843 ldsub = -2.30808644980433e-7   voffl = 0.0   minv = 0.0   pclm = 1.57294391828857 lpclm = -2.18785516397432e-7   pdiblc1 = 1.07192767549886 lpdiblc1 = -2.06957897661431e-7   pdiblc2 = 0.0201843356566257 lpdiblc2 = -3.75248807004432e-9   pdiblcb = -0.538021940443525 lpdiblcb = 1.24906903871122e-7   drout = -0.787931678836857 ldrout = 4.15234616888108e-7   pscbe1 = 800000000.0   pscbe2 = 8.39560530674999e-09 lpscbe2 = 2.51135943258058e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.0571669129457 lbeta0 = -3.4291025292725e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.00654021112577e-08 lagidl = -2.26758158669706e-15   bgidl = 1000000000.0   cgidl = -732.900344667757 lcgidl = 0.000239883874746674 pcgidl = -5.16987882845642e-26   egidl = 5.56577277461714 legidl = -1.26938746649541e-6   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.322483916714286 lkt1 = -6.3986681730524e-8   kt2 = 0.141880867971429 lkt2 = -6.12751947002884e-8   at = 16037.5965142858 lat = 0.0121415255037327   ute = -0.3   ua1 = 4.25248233285714e-10 lua1 = -6.74963727829741e-17   ub1 = 3.927e-19   uc1 = 6.0045e-13   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.35 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.913721522121076+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.66324256720344e-08 wvth0 = 1.69155993604289e-07 pvth0 = -3.9285295422641e-14   k1 = 1.10347180508922 lk1 = -1.52816602548363e-08 wk1 = -5.72768040572178e-06 pk1 = 1.33021368046604e-12   k2 = -0.283048330138908 lk2 = 2.04134281668107e-08 wk2 = 2.48438846261025e-06 pk2 = -5.76981829721993e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 962918.1542418 lvsat = -0.204199461328579 wvsat = -1.86310057530505 pvsat = 4.32692066910572e-7   ua = -2.57310258543751e-09 lua = 8.39493150896677e-17 wua = 5.92992143472816e-15 pua = -1.37718274376557e-21   ub = 7.76621505270878e-18 lub = -1.31806417752505e-24 wub = -2.21435964995498e-23 pub = 5.14269528184495e-30   uc = -5.91444756871381e-13 luc = 1.9596389988357e-19 wuc = 3.57795926866618e-18 puc = -8.3095599443284e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0117342355300624 lu0 = -1.86194218634828e-09 wu0 = -1.53048096805406e-08 pu0 = 3.55443491463779e-15   a0 = -2.49043711907807 la0 = 7.85287231686048e-07 wa0 = 1.07563311679691e-05 pa0 = -2.49808261944264e-12   keta = -0.606361830328397 lketa = 1.46372769792221e-07 wketa = 2.04446480081701e-06 pketa = -4.74812638736145e-13   a1 = 0.0   a2 = -1.53677292901034 la2 = 5.12943445981837e-7   ags = -14.2629578822037 lags = 3.60277587743664e-06 wags = 4.5613559837445e-05 pags = -1.05934299773278e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.213707340242167+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -8.54383439037777e-09 wvoff = 1.10369785769668e-06 pvoff = -2.56326101565051e-13   nfactor = {6.09322934269254+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.83205650742344e-07 wnfactor = -1.20470760156286e-05 pnfactor = 2.79784907509763e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -1.47129769755946 leta0 = 3.83969690020211e-07 weta0 = 1.91274851328237e-06 peta0 = -4.44222452970237e-13   etab = -0.331199875050948 letab = 5.87216957071213e-08 wetab = -5.34318706300601e-07 petab = 1.2409177930737e-13   dsub = 0.354529798969879 ldsub = -1.92353009600516e-08 wdsub = -1.14978382737744e-08 pdsub = 2.67029245421632e-15   voffl = 0.0   minv = 0.0   pclm = 3.10296433617254 lpclm = -5.7412204830806e-07 wpclm = -3.55212547916546e-06 ppclm = 8.24956277657823e-13   pdiblc1 = 1.268202099315 lpdiblc1 = -2.52541258671764e-7   pdiblc2 = 0.0282739368619133 lpdiblc2 = -5.63124132276394e-9   pdiblcb = -0.327552303249288 lpdiblcb = 7.60268039202212e-08 wpdiblcb = 9.59679988184663e-07 ppdiblcb = -2.22878959495971e-13   drout = 1.0   pscbe1 = 556740731.078392 lpscbe1 = 56.4952623921599 wpscbe1 = 715.267926544024 ppscbe1 = -0.000166115969064365   pscbe2 = 5.52404373681349e-09 lpscbe2 = 9.18036016944818e-16 wpscbe2 = 1.00036654589645e-14 ppscbe2 = -2.32328127718631e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 17.4857783887977 lbeta0 = -2.06815326791355e-06 wbeta0 = -2.43048085517142e-06 pbeta0 = 5.64462165247577e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.11679190465832e-09 lagidl = 3.29404698141323e-16 wagidl = 4.76478164317449e-15 pagidl = -1.10658718315577e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.137152910459088 lkt1 = -1.0702851061625e-07 wkt1 = 5.67699514688327e-07 pkt1 = -1.31844238389761e-13   kt2 = -0.0963217202010056 lkt2 = -5.95431101535776e-09 wkt2 = -7.5385572411187e-08 pkt2 = 1.75077714934914e-14   at = 114276.010567883 lat = -0.010673658491317 wat = 0.465813605853004 pat = -1.08181949264119e-7   ute = 0.845481715305048 lute = -2.6603011000759e-07 wute = -3.36811968165697e-06 pute = 7.8222221922706e-13   ua1 = 1.40637147299764e-10 lua1 = -1.397440340339e-18 wua1 = -1.76925323005843e-17 pua1 = 4.10896677908466e-24   ub1 = 2.74580782354632e-19 lub1 = 2.74323614636127e-26 wub1 = 3.47312101465828e-25 pub1 = -8.06608043807281e-32   uc1 = -6.63947539638478e-10 luc1 = 1.54336618757609e-16 wuc1 = 1.21296155250135e-15 puc1 = -2.81701829837571e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.36 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.058106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020121864   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.9074547e-10   ub = 6.7508962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111103   a0 = 1.169205   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.13690013   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22832658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.718041+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.37 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.058106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020121864   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.9074547e-10   ub = 6.7508962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111103   a0 = 1.169205   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.13690013   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22832658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.718041+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.38 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06213291648125+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.24257100477347e-8   k1 = 0.390192585249267 lk1 = 2.64410333808604e-7   k2 = 0.0334579811031172 lk2 = -1.07385655590756e-07 wk2 = 5.29395592033938e-23   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 77362.3059087987 lvsat = -0.192644324783984   ua = -9.54963130039219e-11 lua = -7.66969357677567e-16   ub = 5.39652069525019e-19 lub = 1.09057606774931e-24   uc = -1.12154474749911e-10 luc = 1.09079281016842e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01103391521945 lu0 = 6.15068814490435e-10   a0 = 1.1926370951475 la0 = -1.88680924126788e-7   keta = 0.00982629744199512 lketa = -7.9083709092642e-08 wketa = 4.74336382510877e-24 pketa = -1.952430740422e-29   a1 = 0.0   a2 = 0.8   ags = -0.0316340240020125 lags = 1.35707796182363e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.227296672049727+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -8.29306908322664e-9   nfactor = {1.75682755040487+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.12318728991801e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.118621319005712 lpclm = 2.15310752635537e-6   pdiblc1 = 0.39   pdiblc2 = 0.0001684781660675 lpdiblc2 = 1.88517775900135e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 713696623.183008 lpscbe1 = 349.722254583015   pscbe2 = 1.02399768933739e-08 lpscbe2 = -2.95304653026838e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.1113753017793e-11 lalpha0 = -2.65556694823196e-17   alpha1 = -8.96841316424274e-13 lalpha1 = 7.22209195873408e-18 walpha1 = -6.86488700880216e-34 palpha1 = -1.10489581315083e-39   beta0 = 16.4466505479362 lbeta0 = -5.44890955563207e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37945359045825e-11 lagidl = 2.91535194824076e-16   bgidl = 1709685443.33537 lbgidl = -2875.81786995767   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.435661274676058 lkt1 = -6.97245760515383e-8   kt2 = -0.0539177913697827 lkt2 = 1.00908564946194e-8   at = 134248.740964903 lat = -0.356301614693449 wat = -2.22044604925031e-16   ute = -0.18709643648423 lute = 1.27667076618716e-7   ua1 = 2.03745022542645e-09 lua1 = 5.83086867619045e-16   ub1 = -5.5134482266655e-19 lub1 = -1.50680928618932e-24   uc1 = 3.54684059921587e-10 luc1 = -1.9654421999395e-15 wuc1 = 3.94430452610506e-31 puc1 = -1.50463276905253e-36   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.39 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0617930492405+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.10484854004685e-8   k1 = 0.396175167497855 lk1 = 2.40167456769838e-7   k2 = 0.0288872973925625 lk2 = -8.88641345194465e-08 pk2 = -5.04870979341448e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 35166.4189627955 lvsat = -0.0216563372782503   ua = 2.39821967327358e-10 lua = -2.12576051192203e-15   ub = 5.27340487637494e-19 lub = 1.14046558927195e-24   uc = -1.06505251716063e-10 luc = 8.61872565224953e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01351263572555 lu0 = -9.42930900530992e-9   a0 = 1.269299878692 la0 = -4.99337152105503e-7   keta = 0.0027231515263313 lketa = -5.03000357779148e-08 pketa = 5.04870979341448e-29   a1 = 0.0   a2 = 0.8   ags = 0.084747090339945 lags = 8.8547340589923e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.242704245700565+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.41421633903642e-8   nfactor = {1.7536738301684+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.99539088239589e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.409570498982406 lpclm = 1.27459292557421e-8   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -0.0492804311967633 lpdiblcb = 9.83902073540654e-8   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.00016842862569e-08 lpscbe2 = -1.9874269811267e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.2249091881834e-11 lalpha0 = 1.4916111522228e-16 palpha0 = -9.4039548065783e-38   alpha1 = -1.00818213493928e-10 lalpha1 = 4.1212777291542e-16 walpha1 = -4.62223186652937e-32 palpha1 = 2.057115113939e-37   beta0 = -0.608633512779299 lbeta0 = 1.46230598917253e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.11959196440775e-10 lagidl = 9.63602863189145e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.430536915819335 lkt1 = -9.04897233581801e-8   kt2 = -0.0465295136580214 lkt2 = -1.98482401449209e-8   at = 65916.269111195 lat = -0.0794018339515661   ute = 0.759205248425275 lute = -3.70697730194403e-06 pute = 3.23117426778526e-27   ua1 = 4.6001291289309e-09 lua1 = -9.80151078035454e-15   ub1 = -2.50124286704804e-18 lub1 = 6.39465141486927e-24 pub1 = 5.60519385729927e-45   uc1 = -2.74455005969835e-10 luc1 = 5.83982175845552e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.40 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.067025954293+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.17876781641285e-8   k1 = 0.5473179077703 lk1 = -7.0014173955104e-8   k2 = -0.0306361297303179 lk2 = 3.32924021294949e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -23372.5686226541 lvsat = 0.0984798902210754   ua = -2.24435517749833e-10 lua = -1.17299133797476e-15   ub = 8.0555432378014e-19 lub = 5.69503191545061e-25   uc = -1.00717959024594e-10 luc = 7.43103256074759e-17 wuc = -1.97215226305253e-31   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0114670586675 lu0 = -5.2312878069662e-9   a0 = 0.875203734828998 la0 = 3.09443900464329e-7   keta = -0.0363866141112533 lketa = 2.99627069834588e-8   a1 = 0.0   a2 = 0.8   ags = 0.47871484501648 lags = 7.69558391385948e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21160727277401+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.67638161934739e-9   nfactor = {1.8264322366809+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.4885701869602e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.35141963 leta0 = 8.85377915730091e-07 peta0 = -2.01948391736579e-28   etab = 23.819681025454 letab = -4.90274306567208e-05 wetab = -1.14349447879331e-20 petab = -2.03967875653945e-26   dsub = 0.875672900000001 ldsub = -6.478374993147e-7   voffl = 0.0   minv = 0.0   pclm = 0.19352212829884 lpclm = 4.56129685652495e-7   pdiblc1 = 0.404624957098121 lpdiblc1 = -3.00139658299172e-8   pdiblc2 = -1.12322450000002e-05 lpdiblc2 = 4.64283541175535e-10   pdiblcb = -0.00192751819088942 lpdiblcb = 1.21052310815198e-9   drout = 0.35017133948588 ldrout = 4.30619399739479e-7   pscbe1 = 800000000.0   pscbe2 = 1.07861123141011e-08 lpscbe2 = -3.59726391027389e-15   pvag = 0.0   delta = 0.01   alpha0 = -1.72372784857099e-12 lalpha0 = 1.07038080562564e-16   alpha1 = 1.0e-10   beta0 = 4.0331472627167 lbeta0 = 5.09699778767911e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.2090346350012e-10 lagidl = -1.27219823143757e-16 wagidl = 3.94430452610506e-31   bgidl = 791211102.883898 lbgidl = 428.485552584238   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.500978164719999 lkt1 = 5.40728366094666e-8   kt2 = -0.0625207714580001 lkt2 = 1.29697067362802e-8   at = -12303.6127810001 lat = 0.0811243711225179   ute = -1.72079858075 lute = 1.38259319645412e-6   ua1 = -6.26272093720001e-10 lua1 = 9.24334544022214e-16 wua1 = 3.94430452610506e-31   ub1 = 7.2219766731e-19 lub1 = -2.20631857683278e-25   uc1 = -7.86610627510001e-11 luc1 = 1.82165426432301e-16 puc1 = -9.4039548065783e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.41 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.053353466422+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.74008985092841e-8   k1 = 0.51401774048586 lk1 = -3.49743060312232e-8   k2 = -0.014020275351072 lk2 = 1.58084856699141e-08 wk2 = 9.92616735063633e-24 pk2 = -3.15544362088405e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 88998.418987736 lvsat = -0.0197616948950443   ua = -1.4981191443158e-09 lua = 1.67233342293891e-16   ub = 1.4704150546063e-18 lub = -1.30091858441648e-25   uc = -5.54344501838022e-11 luc = 2.66610704143146e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00614440599032001 lu0 = 3.69436214027711e-10   a0 = 1.350622929424 la0 = -1.90812619113897e-7   keta = -0.00295777191431541 lketa = -5.21255821637371e-9   a1 = 0.0   a2 = 0.75450389119454 la2 = 4.78729620177834e-8   ags = 0.054029874362139 lags = 5.2382762671483e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.231460813028959+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.1214367139142e-8   nfactor = {1.1136174798474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.01197319478732e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -47.9261614871143 letab = 2.64666299062316e-5   dsub = 0.22760894893034 ldsub = 3.40832567506921e-8   voffl = 0.0   minv = 0.0   pclm = 0.63160281715444 lpclm = -4.83765263099056e-9   pdiblc1 = 0.5826111596911 lpdiblc1 = -2.17298701604962e-7   pdiblc2 = 0.00025613852915488 lpdiblc2 = 1.82944515666481e-10   pdiblcb = 0.246873961168832 lpdiblcb = -2.60589091937759e-07 wpdiblcb = -4.30133918527574e-23 ppdiblcb = 1.26217744835362e-29   drout = 0.49368348102824 ldrout = 2.79609753386521e-7   pscbe1 = 800000000.0   pscbe2 = 5.20729698568598e-09 lpscbe2 = 2.27300546734361e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.31478815201679 lbeta0 = 5.91671133399284e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.87973986291398e-11 lagidl = 1.25003731125722e-16   bgidl = 1417577794.2322 lbgidl = -230.604413820174   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.38456890918 lkt1 = -6.84179876677091e-8   kt2 = -0.044680301402 lkt2 = -5.80280299685535e-9   at = 54756.535718 lat = 0.0105607992854846   ute = -0.50539224092 lute = 1.03690383212384e-7   ua1 = -8.36379234399999e-11 lua1 = 3.53351536784276e-16 pua1 = 3.76158192263132e-37   ub1 = 6.1762288776e-19 lub1 = -1.10593777925245e-25   uc1 = 1.7192864804e-10 luc1 = -8.15158426195537e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.42 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.027823558128+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.33021853632807e-8   k1 = 0.063722299604601 lk1 = 2.13698199127367e-7   k2 = 0.148435560935972 lk2 = -7.3906612728752e-08 wk2 = 5.29395592033938e-23 pk2 = 1.26217744835362e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24830.77092048 lvsat = 0.0156744395765614   ua = -3.59445198490802e-10 lua = -4.61591373570344e-16   ub = 4.84174558059204e-19 lub = 4.14552552093013e-25   uc = -8.030900781986e-12 luc = 4.82792082007394e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00947814772352001 lu0 = -1.47159932193986e-9   a0 = 1.61465159268 la0 = -3.36620600196381e-7   keta = 0.065809139972256 lketa = -4.31886039373496e-08 wketa = 5.29395592033938e-23 pketa = -2.52435489670724e-29   a1 = 0.0   a2 = 0.890992217610922 la2 = -2.75017608273777e-8   ags = 1.121025338429 lags = -6.54131493478464e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.19692696556756+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -7.85670838448397e-9   nfactor = {1.1747338499596+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.6744623189886e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.72830100286768 leta0 = -1.31600060726656e-7   etab = -0.000968718832646105 letab = 2.77676297448353e-10   dsub = 0.0323594607981206 ldsub = 1.41908419825294e-7   voffl = 0.0   minv = 0.0   pclm = 0.349339238499881 lpclm = 1.51040432835941e-7   pdiblc1 = -0.0503220228321597 lpdiblc1 = 1.32234217911231e-7   pdiblc2 = -0.00809476346559456 lpdiblc2 = 4.7946716859529e-09 ppdiblc2 = 3.15544362088405e-30   pdiblcb = -0.3461928541026 lpdiblcb = 6.6927905328182e-8   drout = 1.50062087007432 ldrout = -2.76464371152453e-7   pscbe1 = 800000000.0   pscbe2 = 9.4401995944948e-09 lpscbe2 = -6.4585368052796e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.94662656196522 lbeta0 = -3.09500205625848e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.63997097720492e-09 lagidl = 1.57252849167915e-15 wagidl = 7.88860905221012e-31 pagidl = -1.31655367292096e-36   bgidl = 1000000000.0   cgidl = 589.212096506972 lcgidl = -0.0001597153558113   egidl = -1.4304163768928 legidl = 8.45161731224411e-07 pegidl = -5.04870979341448e-28   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.477353150440001 lkt1 = -1.71785399215627e-8   kt2 = -0.048337964648 lkt2 = -3.78288407289455e-9   at = 95243.744212 lat = -0.0117979781948675   ute = -0.33894417636 lute = 1.17706046955753e-8   ua1 = 9.8452460016e-10 lua1 = -2.36533739736159e-16 wua1 = 1.57772181044202e-30   ub1 = 4.4717324952e-19 lub1 = -1.64641583546733e-26   uc1 = 5.29962718026e-11 luc1 = -1.58362703690832e-17 puc1 = -2.35098870164458e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.43 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.978749102600002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.53022529886854e-9   k1 = -0.114773200682002 lk1 = 2.6764721462049e-7   k2 = 0.232565166926557 lk2 = -9.93341972321644e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53540.3814982858 lvsat = 0.00699716074669365   ua = -8.08506000538573e-10 lua = -3.25865889577021e-16   ub = 1.07580025833286e-18 lub = 2.35737825565201e-25   uc = -2.86156636893698e-11 luc = 6.70439257742381e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00756932292285716 lu0 = -8.94670387713112e-10   a0 = -0.792915753000001 la0 = 3.91049777063978e-7   keta = -0.412110446799685 lketa = 1.01259245727362e-7   a1 = 0.0   a2 = 1.225081562433 la2 = -1.28477926674438e-7   ags = -0.24135482835786 lags = 3.46356719402314e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.131437671832573+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.7650388990828e-8   nfactor = {2.72281576313714+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -2.00450689785661e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.660753149102428 leta0 = -1.11184194761085e-7   etab = 0.25974349550927 letab = -7.85207655018953e-08 wetab = 1.01329625037746e-22 petab = -4.76274771527186e-29   dsub = 1.26552967418843 ldsub = -2.30808644980433e-7   voffl = 0.0   minv = 0.0   pclm = 1.57294391828857 lpclm = -2.18785516397433e-7   pdiblc1 = 1.07192767549886 lpdiblc1 = -2.06957897661431e-7   pdiblc2 = 0.0201843356566257 lpdiblc2 = -3.75248807004433e-9   pdiblcb = -0.538021940443526 lpdiblcb = 1.24906903871122e-7   drout = -0.787931678836854 ldrout = 4.15234616888109e-7   pscbe1 = 800000000.0   pscbe2 = 8.39560530674998e-09 lpscbe2 = 2.51135943258058e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.0571669129457 lbeta0 = -3.4291025292725e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.00654021112577e-08 lagidl = -2.26758158669707e-15   bgidl = 1000000000.0   cgidl = -732.900344667756 lcgidl = 0.000239883874746674 wcgidl = 4.33680868994202e-19 pcgidl = 1.03397576569128e-25   egidl = 5.56577277461714 legidl = -1.26938746649541e-6   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.322483916714285 lkt1 = -6.3986681730524e-8   kt2 = 0.141880867971428 lkt2 = -6.12751947002885e-8   at = 16037.5965142858 lat = 0.0121415255037327   ute = -0.3   ua1 = 4.25248233285713e-10 lua1 = -6.74963727829739e-17   ub1 = 3.927e-19   uc1 = 6.0045e-13   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.44 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.879266475602208+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.46343690407162e-08 wvth0 = 1.023010682903e-07 pvth0 = -2.37587070029453e-14   k1 = -6.6368765153714 lk1 = 1.7823600547339e-06 wk1 = 9.29132148665028e-06 pk1 = -2.15784437602413e-12   k2 = 3.17858371044886 lk2 = -7.83526381835416e-07 wk2 = -4.23239688293473e-06 pk2 = 9.8294454928341e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1632652.5933273 lvsat = 0.398603675799113 wvsat = 3.1732208349963 pvsat = -7.36958326382046e-7   ua = 5.80185830296958e-09 lua = -1.86107672651667e-15 wua = -1.03204523500065e-14 pua = 2.39685281512256e-21   ub = -2.60573512465792e-17 lub = 6.53722233052051e-24 wub = 4.34860347811196e-23 pub = -1.00993271756716e-29   uc = 8.29845130820904e-13 luc = -1.34120727503749e-19 wuc = 8.20156308244704e-19 puc = -1.90475561495675e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.022303235794323 lu0 = 6.04302226644096e-09 wu0 = 5.07398726861676e-08 pu0 = -1.17839802522536e-14   a0 = 11.2033036753453 la0 = -2.39498821163322e-06 wa0 = -1.58143489087201e-05 pa0 = 3.67277183360789e-12   keta = 2.72590751499193 lketa = -6.27523459773009e-07 wketa = -4.42131135436785e-06 pketa = 1.02681861287245e-12   a1 = 0.0   a2 = -1.53677292901034 la2 = 5.12943445981838e-7   ags = 49.7279933818863 lags = -1.12586746169894e-05 wags = -7.85514232279249e-05 pags = 1.8243018184723e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {2.20178294956804+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.6952454576677e-07 wvoff = -3.58320404021519e-06 pvoff = 8.32174055911697e-13   nfactor = {-14.4228671680846+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.78151415121007e-06 wnfactor = 2.77613769844702e-05 pnfactor = -6.44738547500432e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.196713726251339 leta0 = -3.41428707987975e-09 weta0 = -1.32378112253404e-06 peta0 = 3.07438899240673e-13   etab = -1.81288206520682 letab = 4.02832012595492e-07 wetab = 2.34066659106917e-06 petab = -5.43603431109677e-13   dsub = 0.338399560259251 ldsub = -1.5489165931179e-08 wdsub = 1.98005058949164e-08 pdsub = -4.5985288905537e-15   voffl = 0.0   minv = 0.0   pclm = -0.630938582369915 lpclm = 2.93050767202995e-07 wpclm = 3.69296126341481e-06 ppclm = -8.57664402699247e-13   pdiblc1 = 1.268202099315 lpdiblc1 = -2.52541258671764e-7   pdiblc2 = 0.0282739368619133 lpdiblc2 = -5.63124132276394e-9   pdiblcb = 1.01960959296333 lpdiblcb = -2.36842116341886e-07 wpdiblcb = -1.65428856088766e-06 ppdiblcb = 3.84196938246234e-13   drout = 1.0   pscbe1 = 1560185215.38 lpscbe1 = -176.547694975498 wpscbe1 = -1231.76778614847 ppscbe1 = 0.00028606944595848   pscbe2 = 1.15029470904632e-08 lpscbe2 = -4.70522434616849e-16 wpscbe2 = -1.59751281687701e-15 ppscbe2 = 3.7101116912997e-22   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 19.379680074625 lbeta0 = -2.50799867713514e-06 wbeta0 = -6.10531715785018e-06 pbeta0 = 1.41791717269059e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.92705945316304e-09 lagidl = -1.30648047275318e-15 wagidl = -8.90277083544718e-15 pagidl = 2.06760620713676e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.155422589333334 lkt1 = -1.74977122414541e-7   kt2 = -0.135173209333333 lkt2 = 3.06867537520108e-9   at = 809579.243136937 lat = -0.172152967132852 wat = -0.883319551129469 pat = 2.05144782512962e-7   ute = -0.890347317 lute = 1.37104031942031e-7   ua1 = 1.14364914775451e-09 lua1 = -2.34339956361952e-16 wua1 = -1.96388907400936e-15 pua1 = 4.56099490215156e-22   ub1 = -5.02711253513174e-20 lub1 = 1.02876943064966e-25 wub1 = 9.77639215257274e-25 pub1 = -2.27049864268995e-31   uc1 = -3.88231150616666e-11 luc1 = 9.15584702061665e-18 wuc1 = -1.84889274661175e-32 puc1 = 2.93873587705572e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.45 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.058106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020121864   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.9074547e-10   ub = 6.7508962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111103   a0 = 1.169205   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.13690013   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22832658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.718041+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.46 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.058106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020121864   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.9074547e-10   ub = 6.7508962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111103   a0 = 1.169205   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.13690013   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22832658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.718041+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.47 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06213291648123+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.24257100477415e-8   k1 = 0.390192585249267 lk1 = 2.64410333808581e-7   k2 = 0.0334579811031168 lk2 = -1.07385655590757e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 77362.3059087992 lvsat = -0.192644324783981   ua = -9.54963130039207e-11 lua = -7.66969357677552e-16   ub = 5.39652069525019e-19 lub = 1.09057606774928e-24   uc = -1.12154474749911e-10 luc = 1.09079281016842e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0110339152194501 lu0 = 6.15068814489588e-10   a0 = 1.1926370951475 la0 = -1.88680924126904e-7   keta = 0.00982629744199499 lketa = -7.90837090926415e-08 wketa = -3.49483808803654e-23 pketa = 3.06866892130974e-28   a1 = 0.0   a2 = 0.8   ags = -0.0316340240020132 lags = 1.35707796182364e-06 pags = 1.29246970711411e-26   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.227296672049725+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -8.29306908321987e-9   nfactor = {1.75682755040486+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.12318728991801e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.118621319005712 lpclm = 2.15310752635535e-6   pdiblc1 = 0.39   pdiblc2 = 0.000168478166067496 lpdiblc2 = 1.88517775900124e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 713696623.182999 lpscbe1 = 349.722254582972   pscbe2 = 1.02399768933738e-08 lpscbe2 = -2.95304653026838e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.11137530177928e-11 lalpha0 = -2.65556694823205e-17   alpha1 = -8.96841316424277e-13 lalpha1 = 7.2220919587341e-18 walpha1 = 2.03576813652807e-33 palpha1 = -1.27880928400003e-38   beta0 = 16.4466505479361 lbeta0 = -5.44890955563202e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37945359045839e-11 lagidl = 2.91535194824068e-16   bgidl = 1709685443.33536 lbgidl = -2875.81786995765   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.435661274676058 lkt1 = -6.97245760515315e-8   kt2 = -0.0539177913697824 lkt2 = 1.00908564946215e-8   at = 134248.740964903 lat = -0.356301614693443 wat = 1.77635683940025e-15   ute = -0.187096436484229 lute = 1.27667076618709e-7   ua1 = 2.03745022542644e-09 lua1 = 5.83086867619158e-16   ub1 = -5.51344822666554e-19 lub1 = -1.50680928618925e-24   uc1 = 3.54684059921588e-10 luc1 = -1.96544219993949e-15 wuc1 = -3.15544362088405e-30   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.48 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06179304924049+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.1048485400455e-8   k1 = 0.396175167497859 lk1 = 2.40167456769843e-7   k2 = 0.0288872973925623 lk2 = -8.88641345194472e-08 wk2 = 2.11758236813575e-22   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 35166.4189627958 lvsat = -0.0216563372782499   ua = 2.39821967327362e-10 lua = -2.12576051192204e-15 pua = -1.20370621524202e-35   ub = 5.27340487637479e-19 lub = 1.14046558927193e-24   uc = -1.06505251716065e-10 luc = 8.61872565224941e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0135126357255499 lu0 = -9.42930900530982e-9   a0 = 1.26929987869201 la0 = -4.99337152105438e-7   keta = 0.00272315152633129 lketa = -5.0300035777915e-8   a1 = 0.0   a2 = 0.8   ags = 0.0847470903399454 lags = 8.85473405899228e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.242704245700562+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.41421633903702e-8   nfactor = {1.75367383016837+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.99539088239589e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.409570498982411 lpclm = 1.27459292557539e-8   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -0.0492804311967636 lpdiblcb = 9.83902073540661e-08 ppdiblcb = -1.61558713389263e-27   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0001684286257e-08 lpscbe2 = -1.98742698112685e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.22490918818339e-11 lalpha0 = 1.49161115222279e-16   alpha1 = -1.00818213493929e-10 lalpha1 = 4.1212777291542e-16 walpha1 = -5.91645678915759e-31 palpha1 = 2.44502824971036e-36   beta0 = -0.608633512779306 lbeta0 = 1.46230598917254e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.11959196440776e-10 lagidl = 9.63602863189145e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.430536915819332 lkt1 = -9.04897233581733e-8   kt2 = -0.0465295136580215 lkt2 = -1.98482401449204e-8   at = 65916.2691111956 lat = -0.0794018339515663   ute = 0.759205248425285 lute = -3.70697730194405e-06 wute = -6.7762635780344e-21 pute = -1.93870456067116e-26   ua1 = 4.60012912893087e-09 lua1 = -9.8015107803546e-15   ub1 = -2.50124286704804e-18 lub1 = 6.39465141486931e-24   uc1 = -2.74455005969834e-10 luc1 = 5.83982175845557e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.49 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.067025954293+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.17876781641437e-8   k1 = 0.547317907770299 lk1 = -7.00141739551048e-8   k2 = -0.0306361297303179 lk2 = 3.3292402129495e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -23372.5686226538 lvsat = 0.0984798902210753 pvsat = -8.470329472543e-22   ua = -2.24435517749834e-10 lua = -1.17299133797476e-15   ub = 8.05554323780143e-19 lub = 5.69503191545091e-25   uc = -1.00717959024593e-10 luc = 7.43103256074759e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0114670586675 lu0 = -5.23128780696602e-9   a0 = 0.875203734829014 la0 = 3.09443900464333e-7   keta = -0.0363866141112532 lketa = 2.99627069834588e-8   a1 = 0.0   a2 = 0.8   ags = 0.478714845016484 lags = 7.69558391385897e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.211607272774014+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.67638161934612e-9   nfactor = {1.82643223668089+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.48857018696007e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.351419630000001 leta0 = 8.85377915730095e-07 weta0 = 1.6940658945086e-21 peta0 = 3.23117426778526e-27   etab = 23.8196810254539 letab = -4.90274306567209e-05 wetab = -2.03287907341032e-20 petab = 1.00166402301343e-25   dsub = 0.875672900000005 ldsub = -6.478374993147e-7   voffl = 0.0   minv = 0.0   pclm = 0.193522128298845 lpclm = 4.56129685652493e-7   pdiblc1 = 0.404624957098122 lpdiblc1 = -3.00139658299147e-8   pdiblc2 = -1.12322449999994e-05 lpdiblc2 = 4.64283541175535e-10   pdiblcb = -0.00192751819088943 lpdiblcb = 1.21052310815196e-9   drout = 0.350171339485883 ldrout = 4.30619399739487e-7   pscbe1 = 800000000.0   pscbe2 = 1.0786112314101e-08 lpscbe2 = -3.59726391027382e-15   pvag = 0.0   delta = 0.01   alpha0 = -1.72372784856996e-12 lalpha0 = 1.07038080562564e-16   alpha1 = 1.0e-10   beta0 = 4.03314726271662 lbeta0 = 5.09699778767909e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.20903463500119e-10 lagidl = -1.2721982314376e-16 wagidl = -3.15544362088405e-30   bgidl = 791211102.883911 lbgidl = 428.485552584243   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.500978164720003 lkt1 = 5.40728366094616e-8   kt2 = -0.0625207714580007 lkt2 = 1.29697067362797e-8   at = -12303.6127809999 lat = 0.0811243711225176   ute = -1.72079858075 lute = 1.38259319645414e-6   ua1 = -6.26272093720003e-10 lua1 = 9.24334544022218e-16   ub1 = 7.22197667309991e-19 lub1 = -2.20631857683285e-25   uc1 = -7.8661062750999e-11 luc1 = 1.82165426432301e-16 puc1 = -1.1284745767894e-36   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.50 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.053353466422+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.74008985092866e-8   k1 = 0.514017740485862 lk1 = -3.49743060312228e-8   k2 = -0.014020275351072 lk2 = 1.58084856699142e-08 wk2 = 7.94093388050907e-23 pk2 = 7.57306469012171e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 88998.4189877352 lvsat = -0.0197616948950445   ua = -1.49811914431579e-09 lua = 1.67233342293891e-16   ub = 1.47041505460631e-18 lub = -1.30091858441637e-25   uc = -5.54344501838019e-11 luc = 2.66610704143146e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00614440599031996 lu0 = 3.69436214027718e-10   a0 = 1.35062292942399 la0 = -1.90812619113909e-7   keta = -0.00295777191431534 lketa = -5.21255821637371e-9   a1 = 0.0   a2 = 0.754503891194531 la2 = 4.78729620177851e-8   ags = 0.0540298743621292 lags = 5.23827626714823e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.23146081302896+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.12143671391422e-8   nfactor = {1.11361747984742+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.01197319478732e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -47.9261614871143 letab = 2.64666299062317e-5   dsub = 0.227608948930339 ldsub = 3.40832567506927e-8   voffl = 0.0   minv = 0.0   pclm = 0.63160281715443 lpclm = -4.83765263099649e-9   pdiblc1 = 0.582611159691091 lpdiblc1 = -2.17298701604966e-7   pdiblc2 = 0.000256138529154876 lpdiblc2 = 1.82944515666479e-10   pdiblcb = 0.24687396116883 lpdiblcb = -2.6058909193776e-07 wpdiblcb = 7.94093388050907e-22 ppdiblcb = -1.0097419586829e-27   drout = 0.493683481028242 ldrout = 2.79609753386524e-7   pscbe1 = 800000000.0   pscbe2 = 5.20729698568606e-09 lpscbe2 = 2.27300546734362e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.31478815201672 lbeta0 = 5.9167113339927e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.87973986291417e-11 lagidl = 1.25003731125722e-16   bgidl = 1417577794.23221 lbgidl = -230.604413820183   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.384568909179997 lkt1 = -6.84179876677052e-8   kt2 = -0.044680301401999 lkt2 = -5.80280299685551e-9   at = 54756.5357179996 lat = 0.0105607992854848   ute = -0.505392240920003 lute = 1.03690383212382e-7   ua1 = -8.36379234400036e-11 lua1 = 3.5335153678428e-16   ub1 = 6.17622887759988e-19 lub1 = -1.10593777925248e-25   uc1 = 1.71928648039997e-10 luc1 = -8.15158426195544e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.51 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.02782355812801+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.33021853632816e-8   k1 = 0.0637222996045992 lk1 = 2.13698199127365e-7   k2 = 0.148435560935972 lk2 = -7.39066127287518e-08 wk2 = -4.2351647362715e-22 pk2 = -1.0097419586829e-28   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24830.7709204806 lvsat = 0.0156744395765613   ua = -3.59445198490799e-10 lua = -4.61591373570348e-16   ub = 4.84174558059189e-19 lub = 4.14552552093007e-25   uc = -8.03090078198605e-12 luc = 4.82792082007406e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00947814772352007 lu0 = -1.47159932193981e-9   a0 = 1.61465159267999 la0 = -3.3662060019638e-07 wa0 = 2.71050543121376e-20   keta = 0.0658091399722567 lketa = -4.31886039373494e-08 pketa = 1.0097419586829e-28   a1 = 0.0   a2 = 0.890992217610929 la2 = -2.75017608273773e-8   ags = 1.12102533842901 lags = -6.54131493478497e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.19692696556756+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -7.85670838448397e-9   nfactor = {1.17473384995958+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.6744623189886e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.728301002867688 leta0 = -1.31600060726652e-7   etab = -0.000968718832646098 letab = 2.77676297448352e-10   dsub = 0.0323594607981192 ldsub = 1.41908419825293e-7   voffl = 0.0   minv = 0.0   pclm = 0.349339238499866 lpclm = 1.51040432835942e-7   pdiblc1 = -0.0503220228321588 lpdiblc1 = 1.32234217911231e-7   pdiblc2 = -0.00809476346559458 lpdiblc2 = 4.79467168595284e-09 wpdiblc2 = 2.64697796016969e-23 ppdiblc2 = -1.26217744835362e-29   pdiblcb = -0.3461928541026 lpdiblcb = 6.69279053281821e-8   drout = 1.50062087007431 ldrout = -2.76464371152454e-7   pscbe1 = 800000000.0   pscbe2 = 9.44019959449483e-09 lpscbe2 = -6.45853680527645e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.9466265619651 lbeta0 = -3.09500205625875e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.63997097720494e-09 lagidl = 1.57252849167913e-15 wagidl = -6.31088724176809e-30 pagidl = 1.05324293833677e-35   bgidl = 1000000000.0   cgidl = 589.21209650697 lcgidl = -0.000159715355811298   egidl = -1.4304163768928 legidl = 8.45161731224408e-07 pegidl = 6.46234853557053e-27   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.477353150440003 lkt1 = -1.71785399215589e-8   kt2 = -0.0483379646479998 lkt2 = -3.78288407289484e-9   at = 95243.7442119997 lat = -0.0117979781948674   ute = -0.338944176360002 lute = 1.1770604695576e-8   ua1 = 9.84524600160006e-10 lua1 = -2.36533739736158e-16   ub1 = 4.47173249520003e-19 lub1 = -1.64641583546722e-26   uc1 = 5.29962718025997e-11 luc1 = -1.58362703690831e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.52 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.978749102600034+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.53022529887701e-9   k1 = -0.114773200682009 lk1 = 2.67647214620489e-7   k2 = 0.232565166926559 lk2 = -9.93341972321644e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53540.3814982846 lvsat = 0.00699716074669432   ua = -8.08506000538553e-10 lua = -3.25865889577027e-16   ub = 1.07580025833284e-18 lub = 2.35737825565195e-25   uc = -2.861566368937e-11 luc = 6.70439257742378e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00756932292285728 lu0 = -8.94670387713082e-10   a0 = -0.792915752999988 la0 = 3.91049777063978e-7   keta = -0.412110446799687 lketa = 1.01259245727362e-07 pketa = -8.07793566946316e-28   a1 = 0.0   a2 = 1.22508156243299 la2 = -1.28477926674435e-7   ags = -0.241354828357856 lags = 3.46356719402314e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.131437671832572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.76503889908293e-8   nfactor = {2.72281576313713+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -2.00450689785654e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.660753149102433 leta0 = -1.11184194761087e-7   etab = 0.259743495509269 letab = -7.85207655018949e-08 wetab = -1.52201232709757e-22 petab = -3.5893171187556e-28   dsub = 1.26552967418841 ldsub = -2.30808644980434e-7   voffl = 0.0   minv = 0.0   pclm = 1.57294391828856 lpclm = -2.18785516397429e-7   pdiblc1 = 1.07192767549886 lpdiblc1 = -2.0695789766143e-7   pdiblc2 = 0.0201843356566256 lpdiblc2 = -3.75248807004427e-9   pdiblcb = -0.538021940443528 lpdiblcb = 1.24906903871123e-7   drout = -0.787931678836856 ldrout = 4.15234616888107e-7   pscbe1 = 800000000.0   pscbe2 = 8.39560530675027e-09 lpscbe2 = 2.51135943258077e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.0571669129454 lbeta0 = -3.4291025292725e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.00654021112577e-08 lagidl = -2.26758158669706e-15   bgidl = 1000000000.0   cgidl = -732.900344667758 lcgidl = 0.000239883874746676 wcgidl = 6.93889390390723e-18   egidl = 5.56577277461713 legidl = -1.2693874664954e-6   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.322483916714276 lkt1 = -6.39866817305236e-8   kt2 = 0.141880867971427 lkt2 = -6.12751947002885e-8   at = 16037.5965142846 lat = 0.0121415255037327   ute = -0.3   ua1 = 4.25248233285717e-10 lua1 = -6.7496372782973e-17   ub1 = 3.927e-19   uc1 = 6.0045e-13   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.53 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.11605232339679+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.64924819287661e-06 wvth0 = -1.1232579137369e-05 pvth0 = 2.60868787659998e-12   k1 = -0.902739525493359 lk1 = 4.50646877793638e-7   k2 = -2.56368768299804 lk2 = 5.50075953392864e-07 wk2 = 5.07210520243404e-06 pk2 = -1.17796092852888e-12   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4559408.87800403 lvsat = -1.03945925648728 wvsat = -6.86009959261064 pvsat = 1.59321010968666e-6   ua = -2.25743347080032e-09 lua = 1.06373728989899e-17 wua = 2.73843880606361e-15 pua = -6.35983243636627e-22   ub = 3.74896168625335e-17 lub = -8.22111618404408e-24 wub = -5.94824347978108e-23 pub = 1.38143791047479e-29   uc = 1.33600441412036e-12 luc = -2.51672677935067e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.129582080334575 lu0 = -2.92312792072824e-08 wu0 = -1.95367833450987e-07 pu0 = 4.53728117441573e-14   a0 = 1.44348176210934 la0 = -1.28337891037547e-7   keta = -0.00270380442853302 lketa = 6.17741888315898e-9   a1 = 0.0   a2 = -1.53677292901034 la2 = 5.12943445981852e-7   ags = 1.25   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {23.2147883423098+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.44964795719326e-06 wvoff = -3.76316735569562e-05 pvoff = 8.7396927618881e-12   nfactor = {-8.07909413784262+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.30821727134753e-06 wnfactor = 1.74822303986169e-05 pnfactor = -4.06012563446596e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.620257499223001 leta0 = 1.86321561237962e-7   etab = -0.368340198895808 letab = 6.73472759378212e-8   dsub = 0.350619438070339 ldsub = -1.83271470136607e-8   voffl = 0.0   minv = 0.0   pclm = 1.64817164034264 lpclm = -2.36256628250438e-7   pdiblc1 = 1.268202099315 lpdiblc1 = -2.52541258671763e-07 wpdiblc1 = -1.35525271560688e-20   pdiblc2 = 0.0282739368619136 lpdiblc2 = -5.631241322764e-9   pdiblcb = -0.00133422461390018 lpdiblcb = 2.64938683702816e-10   drout = 1.0   pscbe1 = 800000000.0   pscbe2 = 1.05170424106796e-08 lpscbe2 = -2.41552974069926e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 15.6117849479665 lbeta0 = -1.63293140923457e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.3271641129399e-10 lagidl = -3.0457761680391e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.155422589333313 lkt1 = -1.74977122414538e-7   kt2 = -0.135173209333331 lkt2 = 3.06867537520087e-9   at = 264438.778533336 lat = -0.0455479102119174   ute = -0.890347316999993 lute = 1.37104031942033e-7   ua1 = -6.83645576666612e-11 lua1 = 4.71417426261802e-17   ub1 = 5.53078699000011e-19 lub1 = -3.72468301918588e-26   uc1 = -3.88231150616666e-11 luc1 = 9.15584702061669e-18 puc1 = -1.17549435082229e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.54 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.19502309645385+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.17746405562987e-7   k1 = 0.211457885045446 wk1 = 3.36473287879396e-7   k2 = 0.0723289084254723 wk2 = -8.30275879575476e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 47898.4761652631 wvsat = 0.00880979391752629   ua = 3.50256721460063e-09 wua = -5.87366795324252e-15   ub = -6.96006155458555e-19 wub = 2.18052518291122e-24   uc = -2.82327878570129e-10 wuc = 2.92179268537876e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0298822227119655 wu0 = -2.98539685832044e-8   a0 = 0.81281766177646 wa0 = 5.66781387395949e-7   keta = -0.0204172261683982 wketa = 3.24784858007115e-8   a1 = 0.0   a2 = 0.8   ags = -0.0941680993956615 wags = 3.67479866969495e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.295394474035831+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.0666157282925e-7   nfactor = {2.42308848610523+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.12127382063192e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.601305931892396 wpclm = -7.19690004029532e-7   pdiblc1 = 0.39   pdiblc2 = -0.000965213633347046 wpdiblc2 = 1.84020230892147e-9   pdiblcb = 0.590565230769231 wpdiblcb = -9.78965518997354e-7   drout = 0.56   pscbe1 = 625221853.746353 wpscbe1 = 209.777675186624   pscbe2 = 7.10710630075385e-09 wpscbe2 = 4.39912840444247e-15   pvag = 0.0   delta = 0.01   alpha0 = 7.26498616043031e-11 walpha0 = -8.72054212064207e-17   alpha1 = 2.57133538660002e-16 walpha1 = -3.08650808824318e-22   beta0 = -52.8626332593476 wbeta0 = 9.9464344130651e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -4.37589193242769e-11 wagidl = 2.28627313616986e-16   bgidl = 2437598871.19 wbgidl = -1725.62496775043   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.132568212224769 wkt1 = -4.95795618647931e-7   kt2 = -0.0532205288042554 wkt2 = 8.84093970551331e-10   at = 336226.092307692 wat = -0.391586207598942   ute = 3.17822860644103 wute = -5.32683729574443e-6   ua1 = 9.39173272468985e-09 wua1 = -1.15807372187035e-14   ub1 = -4.53286100891465e-18 wub1 = 6.03441179089292e-24   uc1 = 4.25775345171415e-10 wuc1 = -5.01243365968048e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.55 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.19502309645385+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.17746405562986e-7   k1 = 0.211457885045446 wk1 = 3.36473287879396e-7   k2 = 0.0723289084254723 wk2 = -8.30275879575476e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 47898.476165263 wvsat = 0.00880979391752629   ua = 3.50256721460063e-09 wua = -5.87366795324252e-15   ub = -6.96006155458555e-19 wub = 2.18052518291122e-24   uc = -2.82327878570129e-10 wuc = 2.92179268537876e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0298822227119655 wu0 = -2.98539685832044e-8   a0 = 0.812817661776462 wa0 = 5.66781387395949e-7   keta = -0.0204172261683982 wketa = 3.24784858007115e-8   a1 = 0.0   a2 = 0.8   ags = -0.0941680993956614 wags = 3.67479866969495e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.295394474035831+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.0666157282925e-7   nfactor = {2.42308848610523+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.12127382063192e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.601305931892396 wpclm = -7.19690004029532e-7   pdiblc1 = 0.39   pdiblc2 = -0.000965213633347047 wpdiblc2 = 1.84020230892147e-9   pdiblcb = 0.590565230769231 wpdiblcb = -9.78965518997354e-7   drout = 0.56   pscbe1 = 625221853.746353 wpscbe1 = 209.777675186624   pscbe2 = 7.10710630075384e-09 wpscbe2 = 4.39912840444247e-15   pvag = 0.0   delta = 0.01   alpha0 = 7.26498616043031e-11 walpha0 = -8.72054212064207e-17   alpha1 = 2.57133538660002e-16 walpha1 = -3.08650808824318e-22   beta0 = -52.8626332593476 wbeta0 = 9.9464344130651e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -4.3758919324277e-11 wagidl = 2.28627313616986e-16   bgidl = 2437598871.19 wbgidl = -1725.62496775043   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.132568212224769 wkt1 = -4.95795618647932e-7   kt2 = -0.0532205288042554 wkt2 = 8.84093970551331e-10   at = 336226.092307692 wat = -0.391586207598942   ute = 3.17822860644103 wute = -5.32683729574443e-6   ua1 = 9.39173272468985e-09 wua1 = -1.15807372187035e-14   ub1 = -4.53286100891465e-18 wub1 = 6.03441179089292e-24   uc1 = 4.25775345171415e-10 wuc1 = -5.01243365968048e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.56 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.2684167122577+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.90983229101238e-07 wvth0 = 3.28063888437422e-07 pvth0 = -8.88303179253301e-13   k1 = -0.0534379707878849 lk1 = 2.13300580086295e-06 wk1 = 7.05528830780909e-07 pk1 = -2.97172491193991e-12   k2 = 0.149501006631892 lk2 = -6.21408487577954e-07 wk2 = -1.84549280944343e-07 pk2 = 8.17477341701071e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 106507.123267271 lvsat = -0.471931068366618 wvsat = -0.0463505244046454 pvsat = 4.44164287087478e-7   ua = 5.65104516610224e-09 lua = -1.73000665456332e-14 wua = -9.13902488368774e-15 pua = 2.62934474856791e-20   ub = -2.33187157251006e-18 lub = 1.31723858533951e-23 wub = 4.56673394146251e-24 pub = -1.92143327725834e-29   uc = -3.86377572712144e-10 luc = 8.37833421307177e-16 wuc = 4.36111307135053e-16 puc = -1.15897575026984e-21   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0364388583879319 lu0 = -5.27956237253502e-08 wu0 = -4.04028072588701e-08 pu0 = 8.49418123842588e-14   a0 = 0.639147244481434 la0 = 1.39843640197099e-06 wa0 = 8.80243801684453e-07 pa0 = -2.52407553121771e-12   keta = 0.00897551095684845 lketa = -2.36677461767608e-07 wketa = 1.35305015838325e-09 pketa = 2.50629571272888e-13   a1 = 0.0   a2 = 0.8   ags = -0.56338948079224 lags = 3.77828458380093e-06 wags = 8.45678460568343e-07 pags = -3.85057127791617e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.312767335960326+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.39890505821481e-07 wvoff = 1.3592845838568e-07 pvoff = -2.35664074353566e-13   nfactor = {3.98874593661678+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.26070542462795e-05 wnfactor = -3.54953631573256e-06 pnfactor = 1.95529596783366e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.376003074107086 lpclm = 7.86952960239629e-06 wpclm = 4.09327640465331e-07 ppclm = -9.09112442476026e-12   pdiblc1 = 0.39   pdiblc2 = 0.000404938208145301 lpdiblc2 = -1.10327955745939e-08 wpdiblc2 = -3.76054748130525e-10 ppdiblc2 = 1.78458403738475e-14   pdiblcb = 0.590565230769231 wpdiblcb = -9.78965518997354e-7   drout = 0.56   pscbe1 = 448160911.458528 lpscbe1 = 1425.73773311055 wpscbe1 = 422.295303319595 ppscbe1 = -0.00171124358351033   pscbe2 = 4.64553483935436e-09 lpscbe2 = 1.9821171569054e-14 wpscbe2 = 8.89713322838244e-15 ppscbe2 = -3.62190278575369e-20   pvag = 0.0   delta = 0.01   alpha0 = 8.60982142618045e-11 lalpha0 = -1.08289403547897e-16 walpha0 = -1.03348180905228e-16 palpha0 = 1.29985423785406e-22   alpha1 = -3.65716297596472e-12 lalpha1 = 2.94504354748078e-17 walpha1 = 4.3898836239578e-18 palpha1 = -3.53508950131436e-23   beta0 = -25.2682028678421 lbeta0 = -0.000222197058958987 wbeta0 = 6.63413089024606e-05 pbeta0 = 2.6671472855495e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.57815353139417e-10 lagidl = 9.18410120792927e-16 wagidl = 3.52437774582881e-16 pagidl = -9.96951917639396e-22   bgidl = 3893973861.83689 lbgidl = -11727.0853238115 wbgidl = -3473.78789179841 pbgidl = 0.0140766326680249   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.165684825145648 lkt1 = -2.40160593239469e-06 wkt1 = -9.5635209281287e-07 pkt1 = 3.70851264519931e-12   kt2 = 0.0219334443026304 lkt2 = -6.0515805387211e-07 wkt2 = -1.20630179524341e-07 pkt2 = 9.78462458149331e-13   at = 657813.074397534 lat = -2.58949652542406 wat = -0.83265168951612 pat = 3.55156643930923e-6   ute = 6.82246588377068 lute = -2.93442841067167e-05 wute = -1.11476728570545e-05 pute = 4.68707824027101e-11   ua1 = 1.58801760153951e-08 lua1 = -5.22465220684781e-14 wua1 = -2.20148094140733e-14 pua1 = 8.40176847966617e-20   ub1 = -8.47749959096549e-18 lub1 = 3.17631884098489e-23 wub1 = 1.26053776733047e-23 pub1 = -5.29110140298893e-29   uc1 = 1.14612232741764e-09 luc1 = -5.80040894536326e-15 wuc1 = -1.25866558987653e-15 puc1 = 6.0989478005115e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.57 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.14947132891115+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.08987632052878e-07 wvth0 = 1.3943934496643e-07 pvth0 = -1.23950693344781e-13   k1 = 0.267503688468913 lk1 = 8.32472208731208e-07 wk1 = 2.04632969750931e-07 pk1 = -9.41973165352214e-13   k2 = 0.0737417141812632 lk2 = -3.14413425059941e-07 wk2 = -7.1334320419627e-08 pk2 = 3.58702810419515e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 45605.3680122647 lvsat = -0.225142356946803 wvsat = -0.0166016055865112 pvsat = 3.23614439049126e-7   ua = 2.8870354139134e-09 lua = -6.09962737539423e-15 wua = -4.2100017286477e-15 pua = 6.31984790883011e-21   ub = 2.7478197353803e-19 lub = 2.60959226799655e-24 wub = 4.01656988526817e-25 pub = -2.33642884558835e-30   uc = -2.3622701763048e-10 luc = 2.29386885531389e-16 wuc = 2.06303295809877e-16 puc = -2.27737845033478e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0309117710781382 lu0 = -3.03985228638498e-08 wu0 = -2.76707531860864e-08 pu0 = 3.33484353921993e-14   a0 = 1.20723274370368 la0 = -9.03584085653898e-07 wa0 = 9.8708604676365e-08 pa0 = 6.42895000111932e-13   keta = -0.0241948569116189 lketa = -1.02263070765186e-07 wketa = 4.28091139389126e-08 pketa = 8.26395270106842e-14   a1 = 0.0   a2 = 0.8   ags = -0.157885307053891 lags = 2.13508313429892e-06 wags = 3.85870966986561e-07 pags = -1.98731958070185e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.349300106176825+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.87930168201898e-07 wvoff = 1.69524961219313e-07 pvoff = -3.71805267785632e-13   nfactor = {0.234376719897961+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.60656213158483e-06 wnfactor = 2.41621750177224e-06 pnfactor = -4.62172446837046e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.171078775383046 leta0 = 1.01743220999452e-06 weta0 = 3.99303682803733e-07 peta0 = -1.61807555351565e-12   etab = 0.149496534780054 letab = -8.89453296586732e-07 wetab = -3.49076796979836e-07 petab = 1.41454400702396e-12   dsub = -0.387467076917154 ldsub = 3.839366830168e-06 wdsub = 1.50680635020276e-06 pdsub = -6.1059454849647e-12   voffl = 0.0   minv = 0.0   pclm = 2.54576721232303 lpclm = -3.97019358839815e-06 wpclm = -3.39730514269403e-06 ppclm = 6.33427662436781e-12   pdiblc1 = 0.39   pdiblc2 = -0.00491655990010227 lpdiblc2 = 1.05312078840656e-08 wpdiblc2 = 8.16098757655942e-09 ppdiblc2 = -1.6748329627081e-14   pdiblcb = 0.491553853408408 lpdiblcb = 4.01218160830755e-07 wpdiblcb = -8.6011699435726e-07 ppdiblcb = -4.8160310203315e-13   drout = 0.56   pscbe1 = 800000124.720995 lpscbe1 = -0.000255957789704553 wpscbe1 = -0.000198350307982764 ppscbe1 = 4.07063032586974e-10   pscbe2 = 1.11239898680097e-08 lpscbe2 = -6.43110247162951e-15 wpscbe2 = -1.78486115101291e-15 ppscbe2 = 7.06700909240721e-21   pvag = 0.0   delta = 0.01   alpha0 = -8.10985461069076e-11 lalpha0 = 5.69232498278894e-16 walpha0 = 9.3591358995645e-17 palpha0 = -6.68061448201129e-22   alpha1 = -4.11128381974791e-10 lalpha1 = 1.68062283036427e-15 walpha1 = 4.9350245912591e-16 palpha1 = -2.0173539053029e-21   beta0 = -180.088723194447 lbeta0 = 0.000405173310790856 wbeta0 = 0.000285436555481438 pbeta0 = -6.21112450727985e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.58953163068166e-10 lagidl = -7.7043718162964e-16 wagidl = -2.33772178212598e-16 pagidl = 1.37851326010641e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.366518233862615 lkt1 = -2.44989811949866e-07 wkt1 = -1.01812251690971e-07 pkt1 = 2.45709555791981e-13   kt2 = -0.16676558729441 lkt2 = 1.59496276023776e-07 wkt2 = 1.91217704226992e-07 pkt2 = -2.85220945846823e-13   at = -52303.2602393612 lat = 0.28806742079396 wat = 0.188010688585622 pat = -5.84405537716908e-7   ute = 0.705662476233424 lute = -4.55751031614773e-06 wute = 8.51518655494087e-08 pute = 1.35264705031149e-12   ua1 = 6.30361852672642e-09 lua1 = -1.34399840209229e-14 wua1 = -2.70914811146077e-15 pua1 = 5.78645392277909e-21   ub1 = -1.5087110935634e-18 lub1 = 3.52396400277074e-24 wub1 = -1.5784750895312e-24 pub1 = 4.5654040413432e-30   uc1 = -4.2490916131034e-10 luc1 = 5.65792407614265e-16 wuc1 = 2.39275096944914e-16 puc1 = 2.89281379241176e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.58 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.16010154242119+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.30803413317369e-07 wvth0 = 1.4802296634596e-07 pvth0 = -1.4156637023557e-13   k1 = 0.787566451363998 lk1 = -2.34822955980891e-07 wk1 = -3.82079799851032e-07 pk1 = 2.62104009074031e-13   k2 = -0.146225454651244 lk2 = 1.37012657406389e-07 wk2 = 1.83827737184509e-07 pk2 = -1.6495173616417e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -339537.670060101 lvsat = 0.565264746935943 wvsat = 0.502813864634267 pvsat = -7.42352323803174e-7   ua = 3.19457329001728e-09 lua = -6.73076982886328e-15 wua = -5.4374281792518e-15 pua = 8.83882525009723e-21   ub = 3.0428842392043e-20 lub = 3.11106427091898e-24 wub = 1.23272251460162e-24 pub = -4.04197725401668e-30   uc = -2.83921125641909e-10 luc = 3.27266784839089e-16 wuc = 2.91357559076814e-16 puc = -4.02289861443207e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0308939416770174 lu0 = -3.03619326002055e-08 wu0 = -3.08955861333286e-08 pu0 = 3.99665762343466e-14   a0 = -1.09944593516444 la0 = 3.83028108630246e-06 wa0 = 3.14038844690334e-06 pa0 = -5.59937116433949e-12   keta = -0.24052129640565 lketa = 3.41691350401362e-07 wketa = 3.24646041083194e-07 pketa = -4.95758333862678e-13   a1 = 0.0   a2 = 0.8   ags = 2.90191432875734 lags = -4.14436924969722e-06 wags = -3.85374063000613e-06 pags = 6.71339364194523e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.178652036359697+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.22811385438142e-08 wvoff = -5.24104327330234e-08 pvoff = 8.36600909052911e-14   nfactor = {3.72284216910606+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.55261666729434e-06 wnfactor = -3.01595970813421e-06 pnfactor = 6.52642318541957e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -1.17709669973054 leta0 = 3.08202545311119e-06 weta0 = 1.31311734433552e-06 peta0 = -3.49344324369862e-12   etab = 97.1130061476914 letab = -0.000199882137155117 wetab = -0.000116562200853465 petab = 2.39912114360078e-10   dsub = 3.74219336151477 ldsub = -4.63569989698085e-06 wdsub = -4.55877712231503e-06 pdsub = 6.34210573742564e-12   voffl = 0.0   minv = 0.0   pclm = -0.233307638525297 lpclm = 1.73314332073138e-06 wpclm = 6.78809658694252e-07 ppclm = -2.0309014439777e-12   pdiblc1 = 0.424504163518837 lpdiblc1 = -7.08109280523882e-08 wpdiblc1 = -3.16149396654409e-08 ppdiblc1 = 6.48815386238235e-14   pdiblc2 = -0.000707535765504331 lpdiblc2 = 1.8932675670059e-09 wpdiblc2 = 1.10736783570181e-09 ppdiblc2 = -2.27258788924419e-15   pdiblcb = 1.33237500564487 lpdiblcb = -1.32435116309846e-06 wpdiblcb = -2.12201095424775e-06 ppdiblcb = 2.10810994389439e-12   drout = 0.841929903710429 ldrout = -5.785886713804e-07 wdrout = -7.82069314483351e-07 pdrout = 1.60499627616326e-12   pscbe1 = 800000000.0   pscbe2 = 1.20216486261499e-08 lpscbe2 = -8.27331637441139e-15 wpscbe2 = -1.96493789204666e-15 ppscbe2 = 7.43657032365653e-21   pvag = 0.0   delta = 0.01   alpha0 = 2.97574274720816e-10 lalpha0 = -2.07896147555055e-16 walpha0 = -4.75989236841829e-16 palpha0 = 5.00856342542157e-22   alpha1 = 7.31663186355178e-10 lalpha1 = -6.64663166199931e-16 walpha1 = -1.00456693807897e-15 palpha1 = 1.05704852862503e-21   beta0 = 26.3241824526263 lbeta0 = -1.84361299330108e-05 wbeta0 = -3.54505968545501e-05 pbeta0 = 3.74259614434802e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -3.44226665395137e-10 lagidl = 4.67434399075375e-16 wagidl = 8.98755943774856e-16 pagidl = -9.45709650545486e-22   bgidl = 148595174.707274 lbgidl = 1747.28959287322 wbgidl = 1021.98565513074 pbgidl = -0.00209736290684248   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.73219955821118 lkt1 = 5.05477126175208e-07 wkt1 = 3.67723451825763e-07 pkt1 = -7.17891805000314e-13   kt2 = -0.174235559221915 lkt2 = 1.74826473622195e-07 wkt2 = 1.77665858492876e-07 pkt2 = -2.57409265301902e-13   at = -22962.9816268098 lat = 0.227854039393302 wat = 0.0169521506945451 pat = -2.33351850739712e-7   ute = -5.22865375863422 lute = 7.62114863664575e-06 wute = 5.57872519942956e-06 pute = -9.92150036913072e-12   ua1 = -2.36422088777952e-09 lua1 = 4.34852874262096e-15 wua1 = 2.7639506881199e-15 pua1 = -5.44567477696876e-21   ub1 = -2.17153118308332e-19 lub1 = 8.7337318895935e-25 wub1 = 1.49389858847984e-24 pub1 = -1.7398533327392e-30   uc1 = -5.57910367762927e-10 luc1 = 8.38743202548142e-16 wuc1 = 7.62175186574189e-16 puc1 = -1.04418991071694e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.59 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.04663136946604+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.14052181165277e-08 wvth0 = -1.06905016825162e-08 pvth0 = 2.54387655031184e-14   k1 = 0.888621216951653 lk1 = -3.41157125687144e-07 wk1 = -5.95751462925023e-07 pk1 = 4.86938520841997e-13   k2 = -0.12508166753965 lk2 = 1.14764255424724e-07 wk2 = 1.76626729402167e-07 pk2 = -1.57374526132255e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 404023.93779126 lvsat = -0.217142749994397 wvsat = -0.501001526885326 pvsat = 3.13905395215577e-7   ua = -5.18117064149463e-09 lua = 2.08254809286261e-15 wua = 5.85734905125165e-15 pua = -3.04602502725942e-21   ub = 4.43113086377523e-18 lub = -1.51954362616734e-24 wub = -4.7085809006866e-24 pub = 2.20971767559644e-30   uc = 1.51614470447134e-11 luc = 1.25592413075996e-17 wuc = -1.12272340468344e-16 puc = 2.24268749438883e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.0040847319788023 lu0 = 6.44413190341522e-09 wu0 = 1.62679320732972e-08 pu0 = -9.66090565394793e-15   a0 = 4.67927866553032 la0 = -2.2503414237064e-06 wa0 = -5.29373497295931e-06 pa0 = 3.27537616534706e-12   keta = 0.119648986342595 lketa = -3.7295308428499e-08 wketa = -1.94987927728745e-07 pketa = 5.10228723819038e-14   a1 = 0.0   a2 = 0.614474777614864 la2 = 1.95217616578202e-07 wa2 = 2.22695608845485e-07 pa2 = -2.34329895538401e-13   ags = -2.23490807860776 lags = 1.26081617069585e-06 wags = 3.64021750916917e-06 pags = -1.17207135229501e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.252615821151638+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.55467362570129e-08 wvoff = 3.36439137089199e-08 pvoff = -6.88999275781804e-15   nfactor = {-2.11890372466687+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.59431955720697e-06 wnfactor = 5.14084720914592e-06 pnfactor = -2.05651979564002e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 3.14566924099326 leta0 = -1.46657474865384e-06 weta0 = -4.22344941988597e-06 peta0 = 2.33237037798609e-12   etab = -195.3892353176 letab = 0.000107901298911046 wetab = 0.000234518223885075 petab = -1.29509805008078e-10   dsub = -1.62006839684928 ldsub = 1.00670250242541e-06 wdsub = 2.93845773175078e-06 pdsub = -1.54680715712114e-12   voffl = 0.0   minv = 0.0   pclm = 2.29887695195659 lpclm = -9.31330189311052e-07 wpclm = -2.65155308828569e-06 ppclm = 1.47344944399272e-12   pdiblc1 = 0.427355348122473 lpdiblc1 = -7.38110670932721e-08 wpdiblc1 = 2.46911421490951e-07 ppdiblc1 = -2.28195875218462e-13   pdiblc2 = 0.00146102414728694 lpdiblc2 = -3.88584421309325e-10 wpdiblc2 = -1.91619249354469e-09 ppdiblc2 = 9.08932302283136e-16   pdiblcb = 1.08365474940402 lpdiblcb = -1.06263701451082e-06 wpdiblcb = -1.33077616748756e-06 ppdiblcb = 1.27553867816949e-12   drout = -0.489833647420856 ldrout = 8.22750202952636e-07 wdrout = 1.5641386289667e-06 pdrout = -8.63784608876459e-13   pscbe1 = 800000000.0   pscbe2 = -1.56536734976649e-09 lpscbe2 = 6.02352607713475e-15 wpscbe2 = 1.07709216257484e-14 ppscbe2 = -5.96464870292669e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.9552904609923 lbeta0 = 1.94465108294209e-06 wbeta0 = 2.16208014381572e-06 pbeta0 = -2.15171463931129e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.61843437099761e-10 lagidl = -4.85971523784164e-16 wagidl = -9.23423430511296e-16 pagidl = 9.71665840791498e-22   bgidl = 2702809650.58545 lbgidl = -940.364709868263 wbgidl = -2043.97131026148 pbgidl = 0.00112876884829273   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.0316374844488032 lkt1 = -2.9826505510446e-07 wkt1 = -6.61914753761633e-07 pkt1 = 3.65537789361586e-13   kt2 = 0.0439310255276992 lkt2 = -5.47377880144932e-08 wkt2 = -1.40923218727566e-07 pkt2 = 7.78238610797674e-14   at = 295596.566586196 lat = -0.107348015296996 wat = -0.383020472939303 pat = 1.8751654267064e-7   ute = 4.85124155167488 lute = -2.98535064435983e-06 wute = -8.51893433664761e-06 pute = 4.91266319408974e-12   ua1 = 3.10726156794236e-09 lua1 = -1.40880037103519e-15 wua1 = -5.07465402609881e-15 pua1 = 2.80244216333489e-21   ub1 = 1.2848140462529e-18 lub1 = -7.07061246180058e-25 wub1 = -1.06106892672974e-24 pub1 = 9.48593350367472e-31   uc1 = 4.76510747364352e-10 luc1 = -2.49719174896732e-16 wuc1 = -4.84392811741102e-16 puc1 = 2.67502539534342e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.60 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08304529307106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.15145525299325e-08 wvth0 = 8.78220076545144e-08 pvth0 = -2.89640781906923e-14   k1 = -1.04243763873834 lk1 = 7.25256609955666e-07 wk1 = 1.75918389149556e-06 pk1 = -8.13558044089289e-13   k2 = 0.56298544934348 lk2 = -2.65215993404166e-07 wk2 = -6.59280327038634e-07 pk2 = 3.04249294437782e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -24509.9827663891 lvsat = 0.0195121078961208 wvsat = 0.0784691761755704 pvsat = -6.10324425488177e-9   ua = 6.24367027787911e-10 lua = -1.12351944623499e-15 wua = -1.56460793844924e-15 pua = 1.05269876660397e-21   ub = -2.36296698699699e-19 lub = 1.05801057321651e-24 wub = 1.14580304822328e-24 pub = -1.0233248795014e-30   uc = 1.15651633756711e-10 luc = -4.29357608727944e-17 wuc = -1.96698790905193e-16 puc = 6.90507912124856e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111233755357085 lu0 = -1.95443901472079e-09 wu0 = -2.61649167061521e-09 pu0 = 7.67885167661485e-16   a0 = 1.88742064844628 la0 = -7.08557376777856e-07 wa0 = -4.33798867929831e-07 pa0 = 5.91510470897258e-13   keta = 0.458047805537481 lketa = -2.2417368753714e-07 wketa = -6.23797624706719e-07 pketa = 2.87830025870111e-13   a1 = 0.0   a2 = 0.143023136789734 la2 = 4.55573485062394e-07 wa2 = 1.18953427321595e-06 pa2 = -7.6825978006634e-13   ags = -2.7837073077736 lags = 1.56388670340808e-06 wags = 6.20990015430013e-06 pags = -2.59116060529007e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.138804191786444+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.73049393785106e-08 wvoff = -9.24356811529008e-08 pvoff = 6.27365809474585e-14   nfactor = {-0.0979645885708642+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 4.78270065871899e-07 wnfactor = 2.02403876165349e-06 pnfactor = -3.35284148171459e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.46175006198159 leta0 = -5.366421694789e-07 weta0 = -1.16644232474974e-06 peta0 = 6.44159608746771e-13   etab = -0.00414033714532487 letab = 1.24790375468285e-09 wetab = 5.04399016112896e-09 petab = -1.54300337111329e-15   dsub = 0.310674023069738 ldsub = -5.95364837779239e-08 wdsub = -4.42618176400706e-07 pdsub = 3.20368345624165e-13   voffl = 0.0   minv = 0.0   pclm = -0.462216134058132 lpclm = 5.93464139788975e-07 wpclm = 1.29065887216946e-06 ppclm = -7.03609515684914e-13   pdiblc1 = 0.458865277468839 lpdiblc1 = -9.1212205005297e-08 wpdiblc1 = -8.09787143245754e-07 ppdiblc1 = 3.5535851026743e-13   pdiblc2 = 0.00455466058453075 lpdiblc2 = -2.09702348832215e-09 wpdiblc2 = -2.01170393668497e-08 ppdiblc2 = 1.09602225821377e-14   pdiblcb = -2.07896974906161 lpdiblcb = 6.83900226395339e-07 wpdiblcb = 2.75572554700723e-06 ppdiblcb = -9.8120328814826e-13   drout = 0.926721425720039 ldrout = 4.04675796960875e-08 wdrout = 9.12702243907607e-07 pdrout = -5.04033425282269e-13   pscbe1 = 799735287.658709 lpscbe1 = 0.146185537491419 wpscbe1 = 0.42098585433996 ppscbe1 = -2.32486491158305e-7   pscbe2 = 9.41899143944953e-09 lpscbe2 = -4.25091736982589e-17 wpscbe2 = 3.37284360341928e-17 ppscbe2 = -3.51089242593589e-23   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 13.7342633643081 lbeta0 = -1.79898925010373e-06 wbeta0 = -6.02367652140699e-06 pbeta0 = 2.3688121787613e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.29656824641027e-08 lagidl = 6.9845099624736e-15 wagidl = 1.64215179797532e-14 pagidl = -8.6069566384372e-21   bgidl = 2032046217.33301 lbgidl = -569.940299198634 wbgidl = -1641.31697223723 pbgidl = 0.000906405808699206   cgidl = 1479.35665114481 lcgidl = -0.000651291455098162 wcgidl = -0.0014156433507863 pcgidl = 7.8177913096828e-10   egidl = -6.14077192796793 legidl = 3.44642261181679e-06 wegidl = 7.49112431343454e-06 pegidl = -4.13692096422403e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.395044505664006 lkt1 = -6.26329128385921e-08 wkt1 = -1.30899734298519e-07 pkt1 = 7.22884619682174e-14   kt2 = 0.112640181387218 lkt2 = -9.26819383738214e-08 wkt2 = -2.5601194869903e-07 pkt2 = 1.41380806585399e-13   at = 194118.615915117 lat = -0.0513075273845472 wat = -0.15724586973777 pat = 6.28340984748153e-8   ute = -0.435543247376216 lute = -6.57607465774578e-08 wute = 1.53626545108596e-07 pute = 1.23302155066042e-13   ua1 = 1.73099554177447e-09 lua1 = -6.48767091946157e-16 wua1 = -1.18715170423264e-15 pua1 = 6.55596218600546e-22   ub1 = -2.92607474568689e-19 lub1 = 1.6405874674302e-25 wub1 = 1.17651190207204e-24 pub1 = -2.87094999272508e-31   uc1 = 5.28916743340352e-11 luc1 = -1.57785071492506e-17 wuc1 = 1.66346814246447e-19 puc1 = -9.18638637399007e-26   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.61 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.943557950508733+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.06445203481323e-08 wvth0 = -5.59663261488754e-08 pvth0 = 1.44949391830467e-14   k1 = 3.3461237359621 lk1 = -6.01155345617919e-07 wk1 = -5.50404505716521e-06 pk1 = 1.38170206304079e-12   k2 = -1.07256388039142 lk2 = 2.29117342662899e-07 wk2 = 2.07561485168605e-06 pk2 = -5.22353629065502e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 281286.121432051 lvsat = -0.0729126240251283 wvsat = -0.362195938544291 pvsat = 1.27084702013393e-7   ua = -7.98045213331323e-09 lua = 1.47722691147371e-15 wua = 1.14059203105397e-14 pua = -2.86755260295519e-21   ub = 7.77722471479015e-18 lub = -1.36402017936091e-24 wub = -1.06576251274607e-23 pub = 2.54417866260184e-30   uc = -1.15086505512107e-10 luc = 2.68032265542311e-17 wuc = 1.37519093528642e-16 puc = -3.19642248324502e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00323185104142708 lu0 = 2.38432773163241e-09 wu0 = 1.71776707766822e-08 pu0 = -5.21476187289701e-15   a0 = -2.92587233668893 la0 = 7.46226734928366e-07 wa0 = 3.39215219537418e-06 pa0 = -5.64856456328936e-13   keta = -1.27106090125727 lketa = 2.98437315330626e-07 wketa = 1.36603374493762e-06 pketa = -3.13582576785303e-13   a1 = 0.0   a2 = 5.04885837403072 la2 = -1.02718087454703e-06 wa2 = -6.08115186463342e-06 pa2 = 1.42925421029567e-12   ags = 6.17467007978096 lags = -1.14372015333857e-06 wags = -1.02037393279134e-05 pags = 2.36974703273258e-12   b0 = 0.0   b1 = 2.15190841520271e-23 lb1 = -6.50399255136111e-30 wb1 = -3.42229228231614e-29 pb1 = 1.03436388628408e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.369564760658885+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 2.24408272392028e-08 wvoff = 3.78705939594524e-07 pvoff = -7.96626759321055e-14   nfactor = {0.161997410715806+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.99698371321501e-07 wnfactor = 4.07260310057366e-06 pnfactor = -9.54448379659708e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -1.65892834541578 leta0 = 4.06561034408104e-07 weta0 = 3.68911056810632e-06 peta0 = -8.23397264248723e-13   etab = 0.737798568669285 letab = -2.22997936955442e-07 wetab = -7.60275937321192e-07 petab = 2.29769587470926e-13   dsub = -0.433213733060409 ldsub = 1.65298383298121e-07 wdsub = 2.70160031495369e-06 pdsub = -6.2994968385826e-13   voffl = 0.0   minv = 0.0   pclm = 4.29900978332007 lpclm = -8.45583065157167e-07 wpclm = -4.33540484579776e-06 ppclm = 9.9682886062465e-13   pdiblc1 = -0.2132435630158 lpdiblc1 = 1.11927987269301e-07 wpdiblc1 = 2.04387490654851e-06 ppdiblc1 = -5.07140868648536e-13   pdiblc2 = -0.0411319423000725 lpdiblc2 = 1.1711432427329e-08 wpdiblc2 = 9.75144775442464e-08 ppdiblc2 = -2.45930799836227e-14   pdiblcb = 0.0302729004910591 lpdiblcb = 4.63964002665916e-08 wpdiblcb = -9.03788950528967e-07 ppdiblcb = 1.24859352130574e-13   drout = 1.261709193857 ldrout = -6.07801283089331e-08 wdrout = -3.2596508710986e-06 pdrout = 7.57031097256553e-13   pscbe1 = 800945401.218897 lpscbe1 = -0.219562815280369 wpscbe1 = -1.5035209083544 ppscbe1 = 3.49182206319659e-7   pscbe2 = 7.71449613059147e-09 lpscbe2 = 4.72662601936903e-16 wpscbe2 = 1.0832034767438e-15 ppscbe2 = -3.52305408988553e-22   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.29481518509999 lbeta0 = 1.47288885924653e-07 wbeta0 = 4.39311214755318e-06 pbeta0 = -7.79589278911226e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.07371773628804e-08 lagidl = -9.24680350021327e-15 wagidl = -4.87789252493237e-14 pagidl = 1.10994209244487e-20   bgidl = -2655720763.45304 lbgidl = 846.904456375084 wbgidl = 5813.88355874322 pbgidl = -0.00134687636538592   cgidl = -3911.98803980289 lcgidl = 0.000978204738327943 wcgidl = 0.00505586910995109 pcgidl = -1.17419020970237e-9   egidl = 22.3884711713141 legidl = -5.1763414102395e-06 wegidl = -2.67540154051234e-05 pegidl = 6.21343279973208e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.02571946897517 lkt1 = 1.27984180097464e-07 wkt1 = 1.11839220765631e-06 pkt1 = -3.05301282444037e-13   kt2 = -0.413026581929816 lkt2 = 6.61971611714089e-08 wkt2 = 8.82498283746834e-07 pkt2 = -2.02725941599737e-13   at = -215136.754568403 lat = 0.0723870435565033 wat = 0.367648637827926 pat = -9.58115921753635e-8   ute = -0.968551602761329 lute = 9.53372977792051e-08 wute = 1.06323251226501e-06 pute = -1.51619881265214e-13   ua1 = -2.07856111759983e-09 lua1 = 5.02644741453108e-16 wua1 = 3.98193870956139e-15 pua1 = -9.06725175335803e-22   ub1 = 2.50196649076922e-19 wub1 = 2.26630517647887e-25   uc1 = 4.45510581964166e-12 luc1 = -1.13889337175476e-18 wuc1 = -6.13026036300992e-18 puc1 = 1.8112415793356e-24   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.62 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.44396787864496+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.0557218259201e-07 wvth0 = 7.90515622992488e-07 pvth0 = -1.82094568131394e-13   k1 = -3.2833689379107 lk1 = 9.38497921440322e-07 wk1 = 3.78603922342267e-06 pk1 = -7.75854980535784e-13   k2 = 1.78281086875653 lk2 = -4.34023455203469e-07 wk2 = -1.84035833164569e-06 pk2 = 3.87103730951011e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -595155.368436044 lvsat = 0.130634776906308 wvsat = 1.33747299675667 pvsat = -2.67651510527708e-7   ua = 5.21844992385124e-09 lua = -1.58812569898835e-15 wua = -9.15084879756416e-15 pua = 1.90661312501818e-21   ub = -4.59099097353191e-18 lub = 1.50841133674208e-24 wub = 7.44055245161296e-24 pub = -1.65899639289496e-30   uc = 3.33591917721631e-12 luc = -6.99552622891468e-19 wuc = -3.18056884330211e-18 puc = 7.12286855797293e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0220324654519768 lu0 = -3.4831329237452e-09 wu0 = -2.43260668132946e-08 pu0 = 4.42419065621197e-15   a0 = -1.07274389444548 la0 = 3.15850626116418e-07 wa0 = 4.00168500859839e-06 pa0 = -7.06416185470565e-13   keta = -1.08190040848 lketa = 2.54506115006555e-07 wketa = 1.71630269348579e-06 pketa = -3.94930088202975e-13   a1 = 0.0   a2 = -4.5029579150946 la2 = 1.1911615958883e-06 wa2 = 4.71727881822609e-06 pa2 = -1.07860572678367e-12   ags = 1.25   b0 = 0.0   b1 = -5.02111963547295e-23 lb1 = 1.01548629843696e-29 wb1 = 7.98534865873761e-29 pb1 = -1.61498086878907e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.02265169278509+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.74115695616988e-07 wvoff = 9.14392525225136e-07 pvoff = -2.04072135638716e-13   nfactor = {5.82072780098981+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.14502150706904e-07 wnfactor = -4.62338200141351e-06 pnfactor = 1.0651332883811e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -3.19485227379609 leta0 = 7.63268615306932e-07 weta0 = 4.09451246385082e-06 peta0 = -9.17549016722114e-13   etab = -1.05578092555624 letab = 1.93548345521977e-07 wetab = 1.09327287201404e-06 petab = -2.00704148655516e-13   dsub = 0.403478209699053 ldsub = -2.90174635641652e-08 wdsub = -8.40640637490308e-08 pdsub = 1.70013684447952e-14   voffl = 0.0   minv = 0.0   pclm = 4.68690855351625 lpclm = -9.35669839243837e-07 wpclm = -4.83266193508683e-06 ppclm = 1.11231333881241e-12   pdiblc1 = 4.49354646387678 lpdiblc1 = -9.81191048946312e-07 wpdiblc1 = -5.12943350593843e-06 ppdiblc1 = 1.15880979699267e-12   pdiblc2 = 0.11514351911859 lpdiblc2 = -2.45824495589256e-08 wpdiblc2 = -1.38153231254988e-07 ppdiblc2 = 3.01390957110378e-14   pdiblcb = -1.3699431580556 lpdiblcb = 3.71586778351644e-07 wpdiblcb = 2.17657022823867e-06 ppdiblcb = -5.90532504623959e-13   drout = 1.0   pscbe1 = 800000000.0   pscbe2 = 9.64335231116767e-09 lpscbe2 = 2.46992559913488e-17 wpscbe2 = 1.38947497187758e-15 ppscbe2 = -4.23434819832912e-22   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 18.8761673341142 lbeta0 = -2.54239908121883e-06 wbeta0 = -5.19151770945098e-06 pbeta0 = 1.44637391296896e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.69783225572913e-09 lagidl = -1.57364687449312e-15 wagidl = -1.15540929664523e-14 pagidl = 2.45421420057778e-21   bgidl = 929629970.281971 lbgidl = 14.2318459202634 wbgidl = 111.913131576126 pbgidl = -2.26336474693509e-5   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 1.11040017147545 lkt1 = -3.68114653559709e-07 wkt1 = -1.51875069871039e-06 pkt1 = 3.07156697559286e-13   kt2 = -0.181873709857249 lkt2 = 1.25135247026596e-08 wkt2 = 7.42702437493099e-08 pkt2 = -1.50206369065919e-14   at = 726117.448644126 lat = -0.146212656360184 wat = -0.734231688703774 pat = 1.60092400499338e-7   ute = -2.88798505369648 lute = 5.41112280724736e-07 wute = 3.17694756935827e-06 pute = -6.42515407269724e-13   ua1 = -6.70279542066052e-11 lua1 = 3.54802449871754e-17 wua1 = -2.12567025323765e-18 pua1 = 1.85458884254855e-23   ub1 = -5.50101491947602e-19 lub1 = 1.85863641165959e-25 wub1 = 1.75444504366994e-24 pub1 = -3.5482422896694e-31   uc1 = -4.69456664027906e-11 luc1 = 1.07985761714996e-17 wuc1 = 1.29177173949694e-17 puc1 = -2.61251791911079e-24   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.63 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.013621+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.003159553   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.3907199e-9   ub = 1.120565e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0050112152   a0 = 1.2849969   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21197527   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20653591+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4889678+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.64 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.013621+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.003159553   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.3907199e-9   ub = 1.120565e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0050112152   a0 = 1.2849969   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21197527   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20653591+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4889678+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.65 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.995110353976001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.4905221987222e-7   k1 = 0.534330211568017 lk1 = -3.4270500463223e-7   k2 = -0.004244936387451 lk2 = 5.96227478386766e-08 pk2 = 2.52435489670724e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 67893.0195028553 lvsat = -0.101902765767199   ua = -1.96257430632239e-09 lua = 4.60471064032861e-15   ub = 1.47262342609327e-18 lub = -2.83485999710056e-24   uc = -2.30581176929812e-11 luc = -1.27696320938344e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00277973129267591 lu0 = 1.79684506723631e-8   a0 = 1.37246851609192 la0 = -7.04342708374888e-7   keta = 0.0101027219190838 lketa = -2.78807675366248e-8   a1 = 0.0   a2 = 0.8   ags = 0.141135791513957 lags = 5.70416694762887e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.199526856719582+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.64386002138693e-8   nfactor = {1.0316669095341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.68229789414782e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.0349967923963257 lpclm = 2.95815466861526e-07 wpclm = 6.61744490042422e-24 ppclm = 6.31088724176809e-29   pdiblc1 = 0.39   pdiblc2 = 9.165120110643e-05 lpdiblc2 = 3.83437455584577e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799970408.137584 lpscbe1 = 0.119832372482051   pscbe2 = 1.20576370776661e-08 lpscbe2 = -1.03524956742243e-14   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.35796617233013e-10 lagidl = 8.78606223712162e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.631041413047501 lkt1 = 6.87914497691842e-7   kt2 = -0.0785622098265 lkt2 = 2.09988082527966e-07 wkt2 = 5.29395592033938e-23   at = -35859.740561375 lat = 0.369273774917148 wat = -1.38777878078145e-17 pat = -5.29395592033938e-23   ute = -2.464535762125 lute = 9.7032407803207e-6   ua1 = -2.4601156207375e-09 lua1 = 1.77476719661242e-14 wua1 = 3.94430452610506e-31 pua1 = -4.51389830715758e-36   ub1 = 2.02389964278e-18 lub1 = -1.23163859266578e-23   uc1 = 9.7542094152325e-11 luc1 = -7.194437082341e-16 wuc1 = -1.23259516440783e-32 puc1 = -1.88079096131566e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.66 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0333059693055+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.72569497742862e-9   k1 = 0.437981128132815 lk1 = 4.77248942744872e-8   k2 = 0.01431388923153 lk2 = -1.55821233640598e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 31774.755974805 lvsat = 0.0444572147864982   ua = -6.20269965830725e-10 lua = -8.34632727298355e-16   ub = 6.09397920863171e-19 lub = 6.63139513889589e-25   uc = -6.43580479981695e-11 luc = 3.96610325413436e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.007859575909015 lu0 = -2.61631411528468e-9   a0 = 1.2894657788715 la0 = -3.67995447492582e-7   keta = 0.0114689373805169 lketa = -3.34170045767091e-08 wketa = -3.30872245021211e-24   a1 = 0.0   a2 = 0.8   ags = 0.163579482185935 lags = 4.794694063432e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.208070755975015+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.18166442633376e-8   nfactor = {2.2473005115753+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.24374486028843e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.16157665925 leta0 = -3.30568446409198e-7   etab = -0.141315442721079 letab = 2.88987503558393e-7   dsub = 0.86783645 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = -0.284489726177214 lpclm = 1.3068214613246e-06 ppclm = -3.02922587604869e-28   pdiblc1 = 0.39   pdiblc2 = 0.00188226762448545 lpdiblc2 = -3.4216383114769e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799999959.47757 lpscbe1 = 8.31618726806482e-5   pscbe2 = 9.63704199469976e-09 lpscbe2 = -5.43656193439487e-16   pvag = 0.0   delta = 0.01   alpha0 = -3.1286311139205e-12 lalpha0 = 1.26779735309665e-17   alpha1 = 3.00023612205075e-15 lalpha1 = -1.21576858239273e-20   beta0 = 57.7052805 lbeta0 = -0.000112268528969162   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.42001745597948e-11 lagidl = 3.77986806018663e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.451336882665 lkt1 = -4.02919276189324e-8   kt2 = -0.00746425537950002 lkt2 = -7.81181056942088e-8   at = 104326.3427935 lat = -0.198794300055061   ute = 0.776601543575 lute = -3.43063517874099e-06 wute = 1.05879118406788e-22 pute = 6.05845175209737e-28   ua1 = 4.046657518565e-09 lua1 = -8.61935394020239e-15   ub1 = -2.823721046085e-18 lub1 = 7.32735107645062e-24   uc1 = -2.25571752719e-10 luc1 = 5.89892115953299e-16 wuc1 = -9.86076131526265e-32 puc1 = -1.88079096131566e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.67 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.036785263794+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.28660527363897e-8   k1 = 0.46926004108622 lk1 = -1.64670358817483e-8   k2 = 0.006919378327368 lk2 = -4.06790122569682e-10   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 79350.939994737 lvsat = -0.053180675835119   ua = -1.33528734526277e-09 lua = 6.32756684519405e-16   ub = 1.05739618964364e-18 lub = -2.56261797227252e-25   uc = -4.1194400038529e-11 luc = -7.87640183829312e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00515517422749 lu0 = 2.93377530481325e-9   a0 = 1.516776575948 la0 = -8.34492439617252e-7   keta = 0.0299376914507431 lketa = -7.13193758360523e-08 wketa = -6.61744490042422e-24 pketa = -1.26217744835362e-29   a1 = 0.0   a2 = 0.8   ags = -0.30859391207909 lags = 1.44848394950984e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.2223145820134+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.41514801715583e-9   nfactor = {1.2102798493684+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.84473534581047e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.0831533185000001 leta0 = 1.71676937318396e-07 weta0 = -1.65436122510606e-24 peta0 = 3.70764625453876e-29   etab = 0.00633957644215793 letab = -1.40364759342256e-08 petab = -3.15544362088405e-30   dsub = -0.0556729000000002 ldsub = 6.47837499314701e-7   voffl = 0.0   minv = 0.0   pclm = 0.33220110023842 lpclm = 4.1222029648894e-8   pdiblc1 = 0.39816611068281 lpdiblc1 = -1.67588434860219e-8   pdiblc2 = 0.000215   pdiblcb = -0.4354486 lpdiblcb = 4.318916662098e-7   drout = 0.1903966999696 ldrout = 7.58515785264287e-7   pscbe1 = 800000000.0   pscbe2 = 1.0384680832825e-08 lpscbe2 = -2.07799276551018e-15   pvag = 0.0   delta = 0.01   alpha0 = -9.89670377721591e-11 lalpha0 = 2.0936167272649e-16 walpha0 = 1.54074395550979e-32 palpha0 = 2.93873587705572e-38   alpha1 = -1.05230300472244e-10 lalpha1 = 2.15952147059816e-16 walpha1 = -3.45764610328271e-33 palpha1 = 8.15556603068061e-38   beta0 = -3.2093135117666 lbeta0 = 1.27430201893284e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.0451686485778e-10 lagidl = -3.20425739428545e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.425853260994609 lkt1 = -9.25905118066385e-8   kt2 = -0.02622411850237 lkt2 = -3.96183079193406e-8   at = -8840.33437832302 lat = 0.0334512210040727 pat = -1.32348898008484e-23   ute = -0.581080155295499 lute = -6.44342416005898e-7   ua1 = -6.16044655995101e-11 lua1 = -1.88202041034665e-16   ub1 = 1.02739709660346e-18 lub1 = -5.76079174054775e-25   uc1 = 7.70492603980321e-11 luc1 = -3.11597398690384e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.68 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0555375069168+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.25979692966547e-8   k1 = 0.39230733263918 lk1 = 6.45059129126914e-8   k2 = 0.0220640863500564 lk2 = -1.63427031264874e-08 pk2 = 6.31088724176809e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -13354.833943674 lvsat = 0.0443683258511564   ua = -3.01478621726061e-10 lua = -4.55061308161036e-16   ub = 5.08464749041079e-19 lub = 3.21347468626707e-25   uc = -7.83713847927621e-11 luc = 3.12428201304553e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00946790038468001 lu0 = -1.60426060500684e-9   a0 = 0.269127234176 la0 = 4.78337846716944e-7   keta = -0.042793276627178 lketa = 5.21127620716367e-9   a1 = 0.0   a2 = 0.8   ags = 0.7977164370712 lags = 2.8437662878889e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22458745272034+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 9.80676030843885e-9   nfactor = {2.16387861967+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.18944096277421e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.37283926 leta0 = 4.7649694146018e-07 weta0 = 1.05879118406788e-22 peta0 = -1.51461293802434e-28   etab = -0.0147244989625 letab = 8.12804996179789e-9   dsub = 0.827927892698719 ldsub = -2.8192524959698e-7   voffl = 0.0   minv = 0.0   pclm = 0.0898977137915802 lpclm = 2.96184071913877e-7   pdiblc1 = 0.63305449333248 lpdiblc1 = -2.63918499910459e-7   pdiblc2 = -0.0001353343994335 lpdiblc2 = 3.68636919463104e-10   pdiblcb = -0.025   drout = 0.813232760060799 ldrout = 1.03140900885744e-7   pscbe1 = 800000000.0   pscbe2 = 7.40776705674219e-09 lpscbe2 = 1.05444391697652e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.7564952605634 lbeta0 = 1.5208166930559e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.074503006143e-10 lagidl = 3.23512426669293e-16 pagidl = 9.4039548065783e-38   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.51979629787078 lkt1 = 6.26039114505296e-9   kt2 = -0.07347053272126 lkt2 = 1.00964007175868e-8   at = -23493.507926354 lat = 0.0488699202977735 pat = -1.32348898008484e-23   ute = -2.245787417529 lute = 1.10733414772847e-6   ua1 = -1.12037597552098e-09 lua1 = 9.25882868879633e-16 pua1 = -3.76158192263132e-37   ub1 = 4.0084938427308e-19 lub1 = 8.32012704108814e-26   uc1 = 7.2968510559936e-11 luc1 = -2.68657994171508e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.69 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0098817601892+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.38490275656453e-9   k1 = 0.423118796694161 lk1 = 4.74904975685769e-8   k2 = 0.0137463784785832 lk2 = -1.17493071784214e-08 pk2 = 3.15544362088405e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 40861.81075852 lvsat = 0.0144275633308827   ua = -6.790903561776e-10 lua = -2.46527871092314e-16   ub = 7.18259012718401e-19 lub = 2.05490055070753e-25   uc = -4.82159302009282e-11 luc = 1.45896814202972e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00894360557268001 lu0 = -1.31472246514352e-9   a0 = 1.52602766068 la0 = -2.15776615516905e-7   keta = -0.0616310226487128 lketa = 1.56142895833341e-8   a1 = 0.0   a2 = 1.13401084291128 la2 = -1.84455149921854e-7   ags = 2.38969109504528 lags = -5.94780232254691e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21581132448708+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 4.96020492451858e-9   nfactor = {1.58823947858+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.98948589915545e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.1754675e-05 letab = -3.7555105736025e-11 petab = -9.24446373305873e-33   dsub = -0.0580662319993199 ldsub = 2.0735880380864e-7   voffl = 0.0   minv = 0.0   pclm = 0.61301734505696 lpclm = 7.29491738498918e-9   pdiblc1 = -0.21575933957752 lpdiblc1 = 2.04832997617258e-07 ppdiblc1 = 5.04870979341448e-29   pdiblc2 = -0.012204620038981 lpdiblc2 = 7.03381542890374e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = -2.76101316827354e-30   pdiblcb = 0.2167944 lpdiblcb = -1.335292648392e-07 wpdiblcb = -5.29395592033938e-23 ppdiblcb = 1.26217744835362e-29   drout = 1.68708346271852 ldrout = -3.79437032702063e-7   pscbe1 = 800086006.26808 lpscbe1 = -0.0474963595033842   pscbe2 = 9.4470902224852e-09 lpscbe2 = -7.17580260428912e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.71600578840079 lbeta0 = 1.74441696881075e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.149006012286e-10 lagidl = -1.85849402417136e-16   bgidl = 664683394.7904 lbgidl = 185.176248010765   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.50409561108 lkt1 = -2.41020323034767e-9   kt2 = -0.100640511312 lkt2 = 2.51008312044728e-8   at = 63118.8395679999 lat = 0.00103885768044898   ute = -0.30755868992 lute = 3.69609005074905e-8   ua1 = 7.41992727239999e-10 lua1 = -1.02597210639199e-16   ub1 = 6.87531439719999e-19 lub1 = -7.51168879352919e-26   uc1 = 5.303025600552e-11 luc1 = -1.58550379072564e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.70 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.990182871218572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.4310514574145e-9   k1 = -1.23923467564843 lk1 = 5.49925198109818e-7   k2 = 0.656607650835871 lk2 = -2.06049626719505e-07 wk2 = -1.58818677610181e-22 pk2 = 1.26217744835362e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -20455.2662575715 lvsat = 0.0329602206394571   ua = 1.52169257933e-09 lua = -9.11699107868937e-16   ub = -1.10152364545e-18 lub = 7.55506625023544e-25   uc = -5.208859142573e-13 luc = 1.74188149960928e-19 puc = 4.59177480789956e-41   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0110786744665714 lu0 = -1.96003209283995e-9   a0 = -0.0999082610000031 la0 = 2.75651135259423e-7   keta = -0.133033458197126 lketa = 3.71951759107931e-08 wketa = -5.29395592033938e-23   a1 = 0.0   a2 = -0.0172812678455738 la2 = 1.63514831509628e-7   ags = -2.32595109449885 lags = 8.30489610039698e-7   b0 = 0.0   b1 = -6.99165030004571e-24 lb1 = 2.11317736163672e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0540690756469995+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.39252575916536e-8   nfactor = {3.55483752928571+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -3.95441904723902e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.41442843112557 leta0 = -2.79402022308686e-7   etab = 0.104421183830743 letab = -3.15794620520552e-08 wetab = 2.54358038360056e-23 petab = -1.09947488665179e-29   dsub = 1.817459290202 ldsub = -3.59505656598053e-7   voffl = 0.0   minv = 0.0   pclm = 0.687232468463856 lpclm = -1.51360841588819e-8   pdiblc1 = 1.489485774714 lpdiblc1 = -3.10565401461553e-7   pdiblc2 = 0.04010627890221 lpdiblc2 = -8.77678759977865e-9   pdiblcb = -0.722663571428571 lpdiblcb = 1.50415330819286e-7   drout = -1.453869509709 ldrout = 5.69894016543347e-7   pscbe1 = 799692834.756857 lpscbe1 = 0.0713369775630781   pscbe2 = 8.61690083876285e-09 lpscbe2 = 1.79160903861501e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.9546678079829 lbeta0 = -5.02178227903467e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 2187760640.37428 lbgidl = -275.163187926244   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.0939994224285723 lkt1 = -1.26358905576921e-7   kt2 = 0.322172873485714 lkt2 = -1.02691554656943e-7   at = 91147.2159428571 lat = -0.00743252288021695   ute = -0.0827844818571428 lute = -3.09755304600516e-8   ua1 = 1.23874751028571e-09 lua1 = -2.52737866531285e-16   ub1 = 4.39e-19   uc1 = -6.51945563285715e-13 luc1 = 3.70031741504164e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.71 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.463653193136309+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.20851780569442e-07 wvth0 = -3.86207266450123e-07 pvth0 = 8.96939341821774e-14   k1 = 4.31294209122039 lk1 = -7.39528990758099e-07 wk1 = -5.3322094322791e-06 pk1 = 1.2383683151808e-12   k2 = -1.5483953277497 lk2 = 3.06046880036144e-07 wk2 = 2.15826235498421e-06 pk2 = -5.01241324108597e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 441333.968939885 lvsat = -0.0742870967105059 wvsat = 0.0933207403609337 pvsat = -2.16730887036443e-8   ua = -6.21769033973112e-09 lua = 8.85718399402574e-16 wua = 4.5765473273355e-15 pua = -1.06287108094238e-21   ub = 4.54321929120739e-18 lub = -5.55445408814581e-25 wub = -3.52371693492944e-24 pub = 8.1835859211882e-31   uc = 2.41059317296337e-12 luc = -5.06627347692463e-19 wuc = -2.06985173837989e-18 puc = 4.80708577276561e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00703301882047969 lu0 = 2.24628189122467e-09 wu0 = 1.0562751177214e-08 pu0 = -2.4531250216497e-15   a0 = -2.29591064781019 la0 = 7.85657317579382e-07 wa0 = 5.46991591196657e-06 pa0 = -1.27034968114285e-12   keta = 0.837721116560906 lketa = -1.88255778794737e-07 wketa = -5.87919227264425e-07 pketa = 1.36540125097572e-13   a1 = 0.0   a2 = 2.49504997233677 la2 = -4.19956512704039e-07 wa2 = -3.68279534506951e-06 pa2 = 8.55303439324979e-13   ags = 1.25   b0 = 0.0   b1 = 1.63138507001067e-23 lb1 = -3.29936210714167e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.02771145115996+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.82196368624604e-07 wvoff = 9.20466017321894e-07 pvoff = -2.13771789260889e-13   nfactor = {1.03779358410874+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.89123932235833e-07 wnfactor = 1.11782360827495e-06 pnfactor = -2.59606708256599e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 3.4263338047155 leta0 = -7.46652961987333e-07 weta0 = -3.85324281209994e-06 peta0 = 8.94888670410528e-13   etab = 0.214124254412559 letab = -5.7057232273188e-08 wetab = -4.31060604552912e-07 petab = 1.00110807983182e-13   dsub = 0.486772600456405 ldsub = -5.04629877114665e-08 wdsub = -1.84046668942277e-07 pdsub = 4.27435505351613e-14   voffl = 0.0   minv = 0.0   pclm = -3.30259341204063 lpclm = 9.11473047807121e-07 wpclm = 4.7575543261737e-06 ppclm = -1.10490868937356e-12   pdiblc1 = -2.7702066704457 lpdiblc1 = 6.78718351079671e-07 wpdiblc1 = 3.58962854910245e-06 ppdiblc1 = -8.33666103129201e-13   pdiblc2 = -0.0541004842143143 lpdiblc2 = 1.31020736866923e-08 wpdiblc2 = 6.4999180482472e-08 ppdiblc2 = -1.50956046727908e-14   pdiblcb = 4.14606429213322 lpdiblcb = -9.80312634397897e-07 wpdiblcb = -4.44458144981188e-06 ppdiblcb = 1.03222292964866e-12   drout = 1.0   pscbe1 = 800000000.0   pscbe2 = 1.56122487141165e-08 lpscbe2 = -1.44545967275425e-15 wpscbe2 = -5.77530295697411e-15 ppscbe2 = 1.34127368463653e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -2.1968453068734 lbeta0 = 2.55216863243009e-06 wbeta0 = 2.01035193747862e-05 pbeta0 = -4.66890165015848e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.07290060660289e-08 lagidl = -2.46851225579275e-15 wagidl = -1.5192569118228e-14 pagidl = 3.52836782972463e-21   bgidl = 1022863549.20667 lbgidl = -4.62399278220346   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.154854058666668 lkt1 = -1.12225842293077e-7   kt2 = -0.12   at = -612951.160978275 lat = 0.156089396471078 wat = 0.873122262807416 pat = -2.02776533681183e-7   ute = -0.241305546333333 lute = 5.83987711709228e-9   ua1 = -1.90744592958187e-09 lua1 = 4.77943536523883e-16 wua1 = 2.20702409540801e-15 pua1 = -5.12565896989843e-22   ub1 = 9.11507062333334e-19 lub1 = -1.09736457677481e-25   uc1 = 6.96162454833922e-13 luc1 = 5.69430910520019e-20 wuc1 = -4.42692566863037e-17 puc1 = 1.02812249805972e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.72 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.013621+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.003159553   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.3907199e-9   ub = 1.120565e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0050112152   a0 = 1.2849969   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21197527   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20653591+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4889678+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.73 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.013621+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.003159553   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.3907199e-9   ub = 1.120565e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0050112152   a0 = 1.2849969   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21197527   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20653591+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4889678+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.74 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.995110353975999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.49052219872227e-7   k1 = 0.534330211568016 lk1 = -3.4270500463223e-7   k2 = -0.004244936387451 lk2 = 5.96227478386766e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 67893.0195028551 lvsat = -0.101902765767199   ua = -1.96257430632238e-09 lua = 4.60471064032861e-15   ub = 1.47262342609327e-18 lub = -2.83485999710055e-24 wub = -1.46936793852786e-39   uc = -2.30581176929812e-11 luc = -1.27696320938343e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0027797312926759 lu0 = 1.79684506723631e-8   a0 = 1.37246851609192 la0 = -7.04342708374895e-7   keta = 0.0101027219190837 lketa = -2.78807675366248e-8   a1 = 0.0   a2 = 0.8   ags = 0.141135791513957 lags = 5.70416694762886e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.199526856719582+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.64386002138693e-8   nfactor = {1.0316669095341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.68229789414782e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.0349967923963257 lpclm = 2.95815466861526e-07 wpclm = 3.30872245021211e-24   pdiblc1 = 0.39   pdiblc2 = 9.165120110643e-05 lpdiblc2 = 3.83437455584578e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799970408.137583 lpscbe1 = 0.119832372467499   pscbe2 = 1.20576370776661e-08 lpscbe2 = -1.03524956742243e-14   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.35796617233012e-10 lagidl = 8.7860622371217e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.6310414130475 lkt1 = 6.87914497691839e-7   kt2 = -0.0785622098264999 lkt2 = 2.09988082527966e-7   at = -35859.740561375 lat = 0.369273774917148 pat = 5.29395592033938e-23   ute = -2.464535762125 lute = 9.7032407803207e-6   ua1 = -2.4601156207375e-09 lua1 = 1.77476719661242e-14 wua1 = 3.94430452610506e-31 pua1 = -4.51389830715758e-36   ub1 = 2.02389964278e-18 lub1 = -1.23163859266578e-23 wub1 = -7.3468396926393e-40 pub1 = 5.60519385729927e-45   uc1 = 9.7542094152325e-11 luc1 = -7.19443708234101e-16 wuc1 = -2.46519032881566e-32 puc1 = 1.88079096131566e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.75 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0333059693055+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.72569497742524e-9   k1 = 0.437981128132815 lk1 = 4.77248942744872e-8   k2 = 0.01431388923153 lk2 = -1.55821233640599e-08 wk2 = -1.32348898008484e-23   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 31774.755974805 lvsat = 0.0444572147864981   ua = -6.20269965830727e-10 lua = -8.34632727298352e-16   ub = 6.09397920863171e-19 lub = 6.63139513889583e-25   uc = -6.43580479981695e-11 luc = 3.96610325413434e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00785957590901501 lu0 = -2.61631411528468e-9   a0 = 1.2894657788715 la0 = -3.67995447492585e-7   keta = 0.0114689373805169 lketa = -3.34170045767091e-8   a1 = 0.0   a2 = 0.8   ags = 0.163579482185935 lags = 4.79469406343201e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.208070755975015+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.18166442633376e-8   nfactor = {2.2473005115753+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.24374486028843e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.16157665925 leta0 = -3.30568446409198e-7   etab = -0.141315442721079 letab = 2.88987503558393e-7   dsub = 0.86783645 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = -0.284489726177214 lpclm = 1.30682146132459e-06 wpclm = 5.29395592033938e-23 ppclm = -1.0097419586829e-28   pdiblc1 = 0.39   pdiblc2 = 0.00188226762448545 lpdiblc2 = -3.4216383114769e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799999959.47757 lpscbe1 = 8.31618744996376e-5   pscbe2 = 9.63704199469976e-09 lpscbe2 = -5.43656193439512e-16   pvag = 0.0   delta = 0.01   alpha0 = -3.1286311139205e-12 lalpha0 = 1.26779735309665e-17   alpha1 = 3.00023612205075e-15 lalpha1 = -1.21576858239273e-20   beta0 = 57.7052805000001 lbeta0 = -0.000112268528969162   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.42001745597955e-11 lagidl = 3.77986806018663e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.451336882665 lkt1 = -4.02919276189324e-8   kt2 = -0.00746425537950007 lkt2 = -7.81181056942089e-8   at = 104326.3427935 lat = -0.198794300055061   ute = 0.776601543575 lute = -3.43063517874099e-06 pute = 1.41363874215605e-27   ua1 = 4.046657518565e-09 lua1 = -8.61935394020239e-15 pua1 = -6.01853107621011e-36   ub1 = -2.823721046085e-18 lub1 = 7.32735107645062e-24 pub1 = -2.80259692864963e-45   uc1 = -2.25571752719e-10 luc1 = 5.89892115953299e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.76 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.036785263794+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.28660527363914e-8   k1 = 0.469260041086221 lk1 = -1.64670358817475e-8   k2 = 0.006919378327368 lk2 = -4.06790122569695e-10   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 79350.939994737 lvsat = -0.0531806758351191   ua = -1.33528734526277e-09 lua = 6.32756684519405e-16   ub = 1.05739618964364e-18 lub = -2.56261797227254e-25   uc = -4.1194400038529e-11 luc = -7.87640183829322e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00515517422749 lu0 = 2.93377530481325e-9   a0 = 1.516776575948 la0 = -8.34492439617252e-7   keta = 0.0299376914507431 lketa = -7.13193758360523e-08 wketa = -6.61744490042422e-24 pketa = -1.89326617253043e-29   a1 = 0.0   a2 = 0.8   ags = -0.308593912079089 lags = 1.44848394950984e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.2223145820134+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.41514801715583e-9   nfactor = {1.2102798493684+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.84473534581047e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.0831533185 leta0 = 1.71676937318396e-07 weta0 = 8.27180612553028e-24 peta0 = -4.57539325028187e-29   etab = 0.00633957644215792 letab = -1.40364759342256e-08 wetab = -1.65436122510606e-24 petab = -4.73316543132607e-30   dsub = -0.0556728999999998 ldsub = 6.478374993147e-7   voffl = 0.0   minv = 0.0   pclm = 0.332201100238421 lpclm = 4.12220296488949e-8   pdiblc1 = 0.398166110682809 lpdiblc1 = -1.67588434860227e-8   pdiblc2 = 0.000215   pdiblcb = -0.4354486 lpdiblcb = 4.318916662098e-7   drout = 0.1903966999696 ldrout = 7.58515785264288e-7   pscbe1 = 800000000.0   pscbe2 = 1.0384680832825e-08 lpscbe2 = -2.07799276551015e-15   pvag = 0.0   delta = 0.01   alpha0 = -9.8967037772159e-11 lalpha0 = 2.0936167272649e-16 walpha0 = -1.23259516440783e-32 palpha0 = 8.22846045575601e-38   alpha1 = -1.05230300472244e-10 lalpha1 = 2.15952147059816e-16 walpha1 = -3.05440452117663e-32 palpha1 = 2.69651975593902e-38   beta0 = -3.2093135117666 lbeta0 = 1.27430201893284e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.04516864857781e-10 lagidl = -3.20425739428545e-16 wagidl = 3.94430452610506e-31   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.425853260994611 lkt1 = -9.25905118066385e-8   kt2 = -0.0262241185023701 lkt2 = -3.96183079193406e-8   at = -8840.33437832299 lat = 0.0334512210040727 pat = 1.32348898008484e-23   ute = -0.581080155295499 lute = -6.44342416005897e-7   ua1 = -6.16044655995103e-11 lua1 = -1.88202041034665e-16   ub1 = 1.02739709660346e-18 lub1 = -5.76079174054775e-25   uc1 = 7.7049260398032e-11 luc1 = -3.11597398690384e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.77 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0555375069168+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.25979692966547e-8   k1 = 0.39230733263918 lk1 = 6.45059129126914e-8   k2 = 0.0220640863500564 lk2 = -1.63427031264874e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -13354.833943674 lvsat = 0.0443683258511564   ua = -3.0147862172606e-10 lua = -4.55061308161036e-16   ub = 5.08464749041079e-19 lub = 3.21347468626706e-25   uc = -7.8371384792762e-11 luc = 3.12428201304553e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00946790038468 lu0 = -1.60426060500683e-9   a0 = 0.269127234176 la0 = 4.78337846716943e-7   keta = -0.042793276627178 lketa = 5.21127620716361e-9   a1 = 0.0   a2 = 0.8   ags = 0.797716437071198 lags = 2.8437662878889e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22458745272034+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 9.80676030843885e-9   nfactor = {2.16387861967+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.18944096277417e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.37283926 leta0 = 4.7649694146018e-07 peta0 = -5.04870979341448e-29   etab = -0.0147244989625 letab = 8.12804996179789e-9   dsub = 0.82792789269872 ldsub = -2.81925249596979e-7   voffl = 0.0   minv = 0.0   pclm = 0.0898977137915802 lpclm = 2.96184071913877e-7   pdiblc1 = 0.633054493332479 lpdiblc1 = -2.63918499910459e-7   pdiblc2 = -0.000135334399433501 lpdiblc2 = 3.68636919463104e-10   pdiblcb = -0.025   drout = 0.813232760060799 ldrout = 1.03140900885744e-7   pscbe1 = 800000000.0   pscbe2 = 7.40776705674221e-09 lpscbe2 = 1.05444391697652e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.75649526056338 lbeta0 = 1.52081669305577e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.074503006143e-10 lagidl = 3.23512426669293e-16 pagidl = 9.4039548065783e-38   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.519796297870779 lkt1 = 6.26039114505296e-9   kt2 = -0.0734705327212599 lkt2 = 1.00964007175868e-8   at = -23493.5079263541 lat = 0.0488699202977735   ute = -2.245787417529 lute = 1.10733414772847e-6   ua1 = -1.12037597552098e-09 lua1 = 9.25882868879632e-16   ub1 = 4.00849384273079e-19 lub1 = 8.32012704108825e-26   uc1 = 7.2968510559936e-11 luc1 = -2.68657994171507e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.78 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0098817601892+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.38490275656453e-9   k1 = 0.42311879669416 lk1 = 4.74904975685769e-8   k2 = 0.0137463784785832 lk2 = -1.17493071784214e-08 pk2 = -3.15544362088405e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 40861.8107585199 lvsat = 0.0144275633308826   ua = -6.79090356177599e-10 lua = -2.46527871092314e-16   ub = 7.18259012718401e-19 lub = 2.05490055070752e-25   uc = -4.82159302009283e-11 luc = 1.45896814202972e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00894360557267999 lu0 = -1.31472246514352e-9   a0 = 1.52602766068 la0 = -2.15776615516904e-7   keta = -0.0616310226487128 lketa = 1.56142895833341e-08 pketa = -1.26217744835362e-29   a1 = 0.0   a2 = 1.13401084291128 la2 = -1.84455149921854e-7   ags = 2.38969109504528 lags = -5.9478023225469e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21581132448708+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 4.96020492451858e-9   nfactor = {1.58823947858+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.98948589915546e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.1754675e-05 letab = -3.7555105736025e-11 petab = 3.08148791101958e-33   dsub = -0.0580662319993204 ldsub = 2.07358803808641e-7   voffl = 0.0   minv = 0.0   pclm = 0.613017345056959 lpclm = 7.29491738498918e-9   pdiblc1 = -0.21575933957752 lpdiblc1 = 2.04832997617258e-07 ppdiblc1 = 1.0097419586829e-28   pdiblc2 = -0.012204620038981 lpdiblc2 = 7.03381542890373e-09 wpdiblc2 = -3.30872245021211e-24 ppdiblc2 = 3.94430452610506e-31   pdiblcb = 0.2167944 lpdiblcb = -1.335292648392e-07 ppdiblcb = -1.26217744835362e-29   drout = 1.68708346271852 ldrout = -3.79437032702064e-7   pscbe1 = 800086006.26808 lpscbe1 = -0.0474963595033842   pscbe2 = 9.4470902224852e-09 lpscbe2 = -7.17580260428912e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.71600578840079 lbeta0 = 1.74441696881072e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.149006012286e-10 lagidl = -1.85849402417136e-16   bgidl = 664683394.7904 lbgidl = 185.176248010765   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.504095611079999 lkt1 = -2.41020323034725e-9   kt2 = -0.100640511312 lkt2 = 2.51008312044728e-8   at = 63118.8395679999 lat = 0.00103885768044898   ute = -0.30755868992 lute = 3.69609005074905e-8   ua1 = 7.41992727239999e-10 lua1 = -1.02597210639199e-16   ub1 = 6.87531439720001e-19 lub1 = -7.51168879352919e-26   uc1 = 5.30302560055201e-11 luc1 = -1.58550379072564e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.79 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.990182871218572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.43105145741535e-9   k1 = -1.23923467564843 lk1 = 5.49925198109817e-7   k2 = 0.656607650835871 lk2 = -2.06049626719505e-07 wk2 = 1.05879118406788e-22 pk2 = -5.04870979341448e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -20455.2662575715 lvsat = 0.0329602206394571   ua = 1.52169257932999e-09 lua = -9.11699107868936e-16   ub = -1.10152364544999e-18 lub = 7.55506625023544e-25   uc = -5.20885914257299e-13 luc = 1.74188149960928e-19 puc = 4.59177480789956e-41   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0110786744665714 lu0 = -1.96003209283995e-9   a0 = -0.0999082609999959 la0 = 2.75651135259423e-7   keta = -0.133033458197126 lketa = 3.71951759107931e-08 wketa = -2.64697796016969e-23 pketa = -6.31088724176809e-30   a1 = 0.0   a2 = -0.0172812678455703 la2 = 1.63514831509629e-7   ags = -2.32595109449886 lags = 8.30489610039698e-07 pags = 4.03896783473158e-28   b0 = 0.0   b1 = -6.99165030004571e-24 lb1 = 2.11317736163672e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0540690756469999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.39252575916539e-8   nfactor = {3.55483752928572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -3.95441904723902e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.41442843112557 leta0 = -2.79402022308686e-7   etab = 0.104421183830743 letab = -3.15794620520552e-08 wetab = -5.1491993131426e-23 petab = -5.27550730366552e-30   dsub = 1.817459290202 ldsub = -3.59505656598053e-7   voffl = 0.0   minv = 0.0   pclm = 0.68723246846386 lpclm = -1.51360841588815e-8   pdiblc1 = 1.489485774714 lpdiblc1 = -3.10565401461553e-7   pdiblc2 = 0.04010627890221 lpdiblc2 = -8.77678759977866e-9   pdiblcb = -0.722663571428572 lpdiblcb = 1.50415330819286e-7   drout = -1.453869509709 ldrout = 5.69894016543347e-7   pscbe1 = 799692834.756855 lpscbe1 = 0.0713369775639876   pscbe2 = 8.61690083876287e-09 lpscbe2 = 1.79160903861495e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.9546678079828 lbeta0 = -5.02178227903467e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 2187760640.37429 lbgidl = -275.163187926244   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.0939994224285723 lkt1 = -1.26358905576921e-7   kt2 = 0.322172873485714 lkt2 = -1.02691554656943e-07 wkt2 = 5.29395592033938e-23 pkt2 = 1.26217744835362e-29   at = 91147.2159428573 lat = -0.00743252288021695   ute = -0.0827844818571428 lute = -3.09755304600517e-8   ua1 = 1.23874751028571e-09 lua1 = -2.52737866531285e-16   ub1 = 4.39e-19   uc1 = -6.51945563285714e-13 luc1 = 3.70031741504164e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.80 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.18483758958428+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 4.6638247214822e-08 wvth0 = 2.9196006735539e-07 pvth0 = -6.78056819228186e-14   k1 = -6.50856918617489 lk1 = 1.77369125283802e-06 wk1 = 4.84382250474435e-06 pk1 = -1.12494386996934e-12   k2 = 2.79478758953283 lk2 = -7.02626950222303e-07 wk2 = -1.92585925628484e-06 pk2 = 4.4726733125736e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 382881.003583798 lvsat = -0.0607118046773119 wvsat = 0.148287114930055 pvsat = -3.44386444327007e-8   ua = -1.02480521229869e-09 lua = -3.20292821247713e-16 wua = -3.0659362659285e-16 pua = 7.12042236208023e-23   ub = 4.22942712638285e-19 lub = 4.01459984622048e-25 wub = 3.50794210336507e-25 pub = -8.14694997911812e-32   uc = -2.34353150034779e-12 luc = 5.97484828811342e-19 wuc = 2.40069985724254e-18 puc = -5.57545736945578e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00513515867209623 lu0 = -5.79692154183644e-10 wu0 = -8.79621297920261e-10 pu0 = 2.04285889092897e-16   a0 = 14.0853953657945 la0 = -3.01878633493821e-06 wa0 = -9.93428123679981e-06 pa0 = 2.30716727727809e-12   keta = 3.40216085573197 lketa = -7.83828957139041e-07 wketa = -2.99939577776136e-06 pketa = 6.96588673614631e-13   a1 = 0.0   a2 = -1.42135001595434 la2 = 4.89599969776652e-7   ags = -20.8147732369886 lags = 5.12438913087795e-06 wags = 2.07486580559034e-05 pags = -4.81873059287716e-12   b0 = 0.0   b1 = 1.63138507001067e-23 lb1 = -3.29936210714167e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.751464286084213+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.18039898265916e-07 wvoff = 6.60696387899149e-07 pvoff = -1.53442111214862e-13   nfactor = {-19.8652291408444+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.04370463894712e-06 wnfactor = 2.07740270143346e-05 pnfactor = -4.82462235589011e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.27766645502983 leta0 = -2.47640010694282e-07 weta0 = -1.83273874275485e-06 peta0 = 4.25640743833615e-13   etab = -1.60919387230462 letab = 3.6639563942999e-07 wetab = 1.28350060720546e-06 petab = -2.98084031519218e-13   dsub = 0.0842886411872144 ldsub = 4.3011094441087e-08 wdsub = 1.94430007621213e-07 pdsub = -4.51550082599737e-14   voffl = 0.0   minv = 0.0   pclm = -3.7804948174572 lpclm = 1.02246230390528e-06 wpclm = 5.20694996414027e-06 ppclm = -1.20927768052183e-12   pdiblc1 = 1.04711682717833 lpdiblc1 = -2.07828309979028e-7   pdiblc2 = 0.01502168137691 lpdiblc2 = -2.95106541671041e-9   pdiblcb = -0.580442914221889 lpdiblcb = 1.17385578727634e-7   drout = 1.0   pscbe1 = -217736826.640068 lpscbe1 = 236.362253829369 wpscbe1 = 957.031063952007 ppscbe1 = -0.000222263765385406   pscbe2 = -9.42410302174487e-09 lpscbe2 = 4.36905776343739e-15 wpscbe2 = 1.77676854778171e-14 ppscbe2 = -4.12642057842464e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 19.4961738773397 lbeta0 = -2.48588322196913e-06 wbeta0 = -2.95558939730691e-07 pbeta0 = 6.86414948398798e-14   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.83940291468841e-08 lagidl = 6.61753881115981e-15 wagidl = 2.15968631149122e-14 pagidl = -5.01572028039655e-21   bgidl = 1022863549.20667 lbgidl = -4.62399278220437   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.154854058666668 lkt1 = -1.12225842293077e-7   kt2 = -0.12   at = 315554.416833333 lat = -0.059549524436624   ute = -0.241305546333333 lute = 5.83987711709228e-9   ua1 = 4.39572661333334e-10 lua1 = -6.71351020860374e-17   ub1 = 9.11507062333334e-19 lub1 = -1.09736457677481e-25   uc1 = -4.63811524983334e-11 luc1 = 1.09903199477204e-17 wuc1 = 6.16297582203915e-33 puc1 = -2.93873587705572e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.81 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.971013282532601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -3.32490260626636e-8   k1 = 0.52979489926727 wk1 = -2.96727981909484e-8   k2 = -0.0252921628241825 wk2 = 2.22023590371756e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 144457.673409517 wvsat = -0.0696229112328507   ua = -2.80098360977231e-09 wua = 1.10050238850098e-15   ub = 2.35374189659135e-18 wub = -9.62312304244233e-25   uc = 4.5504209095516e-11 wuc = -6.58779609820571e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00107727430803591 wu0 = 3.06985942971414e-9   a0 = 1.3838456786411 wa0 = -7.7136861879896e-8   keta = 0.0044135173140715 wketa = 1.73762583980327e-9   a1 = 0.0   a2 = 0.8   ags = 0.14527025553703 wags = 5.20534047872105e-8   b0 = -9.0807708734e-09 wb0 = 7.08619952875361e-15   b1 = -6.5141632689e-09 wb1 = 5.08334163804531e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20462176335635+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.49370854449485e-9   nfactor = {1.5993249627671+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -8.6117454751064e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = -0.00021574359561109 wpdiblc2 = 6.11469887334373e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 828677844.732781 wpscbe1 = -22.3902982093455   pscbe2 = 1.44112221027286e-08 wpscbe2 = -2.83989760436669e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.901761e-10 walpha0 = 2.2643955802242e-16   alpha1 = -2.901761e-10 walpha1 = 2.2643955802242e-16   beta0 = 108.347547 wbeta0 = -6.11386806660534e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.83183150875686e-09 wagidl = 2.3243098116242e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.603645220000001 wkt1 = 4.52879116044837e-8   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.82 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.9710132825326+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -3.32490260626632e-8   k1 = 0.529794899267269 wk1 = -2.96727981909484e-8   k2 = -0.0252921628241825 wk2 = 2.22023590371756e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 144457.673409517 wvsat = -0.0696229112328507   ua = -2.80098360977231e-09 wua = 1.10050238850098e-15   ub = 2.35374189659135e-18 wub = -9.62312304244233e-25   uc = 4.55042090955161e-11 wuc = -6.58779609820571e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00107727430803591 wu0 = 3.06985942971415e-9   a0 = 1.3838456786411 wa0 = -7.71368618798947e-8   keta = 0.0044135173140715 wketa = 1.73762583980327e-9   a1 = 0.0   a2 = 0.8   ags = 0.14527025553703 wags = 5.20534047872106e-8   b0 = -9.0807708734e-09 wb0 = 7.08619952875361e-15   b1 = -6.5141632689e-09 wb1 = 5.08334163804531e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20462176335635+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.49370854449485e-9   nfactor = {1.5993249627671+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -8.6117454751064e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = -0.000215743595611091 wpdiblc2 = 6.11469887334372e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 828677844.73278 wpscbe1 = -22.390298209345   pscbe2 = 1.44112221027286e-08 wpscbe2 = -2.83989760436669e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.901761e-10 walpha0 = 2.2643955802242e-16   alpha1 = -2.901761e-10 walpha1 = 2.2643955802242e-16   beta0 = 108.347547 wbeta0 = -6.11386806660534e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.83183150875686e-09 wagidl = 2.3243098116242e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60364522 wkt1 = 4.52879116044843e-8   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.83 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.87821360232861+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.47245575324824e-07 wvth0 = -9.12206373208945e-08 pvth0 = 4.6680150095281e-13   k1 = 0.648001189738457 lk1 = -9.51825775002578e-07 wk1 = -8.87033978914535e-08 pk1 = 4.75328733224198e-13   k2 = -0.0408320338706751 lk2 = 1.25130817855023e-07 wk2 = 2.85508220126484e-08 pk2 = -5.11193665550098e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 286325.718274476 lvsat = -1.14235597118755 wvsat = -0.170454437038371 pvsat = 8.11919947846824e-7   ua = -4.87625610220897e-09 lua = 1.67105984003156e-14 wua = 2.27369799952004e-15 pua = -9.44685614645896e-21   ub = 3.51408752060122e-18 lub = -9.34338492851412e-24 wub = -1.59306099737029e-24 pub = 5.07894174898343e-30   uc = 9.3644012957973e-11 luc = -3.87633398672842e-16 wuc = -9.10687643981596e-17 puc = 2.02842470471687e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00621367077905429 lu0 = 5.87084615409063e-08 wu0 = 7.01802109215921e-09 pu0 = -3.17915571092916e-14   a0 = 1.71640646439975 la0 = -2.67786025919957e-06 wa0 = -2.68392734625496e-07 pa0 = 1.54003876252465e-12   keta = 0.0274233316478253 lketa = -1.85280616400269e-07 wketa = -1.35161759071649e-08 pketa = 1.22827318340412e-13   a1 = 0.0   a2 = 0.8   ags = -0.133838972544491 lags = 2.24745532805483e-06 wags = 2.14577162077491e-07 pags = -1.30868078697436e-12   b0 = -5.54286290562165e-08 lb0 = 3.73204216617577e-13 wb0 = 4.32538526270025e-14 pb0 = -2.91230731486803e-19   b1 = -1.16419888917294e-08 lb1 = 4.12904979766488e-14 wb1 = 9.08485164403662e-15 pb1 = -3.22211309351735e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.160277438437183+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.57071279920093e-07 wvoff = -3.06283699053912e-08 pvoff = 2.34599373000647e-13   nfactor = {1.14417913717548+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.66494478809936e-06 wnfactor = -8.7799164366851e-08 pnfactor = 1.35415344817452e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 1.02864882530063 lpclm = -8.26891751271944e-06 wpclm = -8.30018197790176e-07 ppclm = 6.68350822302856e-12   pdiblc1 = 0.39   pdiblc2 = -0.00327272598490768 lpdiblc2 = 2.46155650453368e-08 wpdiblc2 = 2.62539913873592e-09 ppdiblc2 = -1.62166477170934e-14   pdiblcb = -0.225   drout = 0.56   pscbe1 = 857730322.680572 lpscbe1 = -233.937612187761 wpscbe1 = -45.073076385434 ppscbe1 = 0.000182647241788963   pscbe2 = 1.96084258782336e-08 lpscbe2 = -4.18491477208839e-14 wpscbe2 = -5.89227465225824e-15 ppscbe2 = 2.45784817172453e-20   pvag = 0.0   delta = 0.01   alpha0 = -5.21579499463169e-10 lalpha0 = 1.8633164035035e-15 walpha0 = 4.07015709880983e-16 palpha0 = -1.45404305477005e-21   alpha1 = -5.84142018656376e-10 lalpha1 = 2.36708501073937e-15 walpha1 = 4.55836509370944e-16 palpha1 = -1.84715999571749e-21   beta0 = 169.098126166786 lbeta0 = -0.000489178425841699 wbeta0 = -0.000108545528770129 pbeta0 = 3.81731460798107e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -6.02915176132311e-09 lagidl = 2.57455996224848e-14 wagidl = 4.8108310300927e-15 pagidl = -2.00220730757644e-20   bgidl = 1945488487.43339 lbgidl = -7613.30305451611 wbgidl = -737.814021243319 pbgidl = 0.00594105778785837   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54700285679068 lkt1 = -4.560980726557e-07 wkt1 = -6.55796722598327e-08 pkt1 = 8.92732726098356e-13   kt2 = -0.17200126630194 lkt2 = 9.6238207095893e-07 wkt2 = 7.29153732865336e-08 pkt2 = -5.87132304138877e-13   at = -13716.7120777503 lat = 0.19097272881108 wat = -0.0172793609918592 pat = 1.39137613591172e-7   ute = -3.32835490454309 lute = 1.66589224231228e-05 wute = 6.74083168188073e-07 pute = -5.42788147246023e-12   ua1 = -7.00156722846351e-09 lua1 = 5.43165438842747e-14 wua1 = 3.54393175328253e-15 pua1 = -2.8536599652847e-20   ub1 = 6.25355689956512e-18 lub1 = -4.63746139650049e-23 wub1 = -3.30062234557823e-24 pub1 = 2.65774131778259e-29   uc1 = 2.02196721446622e-10 luc1 = -1.56214819828221e-15 wuc1 = -8.16674686492846e-17 puc1 = 6.57606302758922e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.84 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.18040117891601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.77291916588435e-07 wvth0 = 1.14786070429023e-07 pvth0 = -3.67987738479837e-13   k1 = 0.328584964280225 lk1 = 3.42526388696963e-07 wk1 = 8.53675371339286e-08 pk1 = -2.30048994735865e-13   k2 = -0.0144863063200404 lk2 = 1.8371527808056e-08 wk2 = 2.24742959590982e-08 pk2 = -2.64958063901932e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -108841.768260888 lvsat = 0.458958709952973 wvsat = 0.109730414043677 pvsat = -3.23457153656448e-7   ua = 7.12027013125757e-10 lua = -5.93448273581769e-15 wua = -1.03966087858204e-15 pua = 3.97967917381808e-21   ub = 6.2032322155371e-19 lub = 2.38285119595106e-24 wub = -8.52558242952402e-27 pub = -1.34198079446238e-30   uc = -2.15553218926974e-11 luc = 7.9182299580443e-17 wuc = -3.34012014824026e-17 puc = -3.0840507680749e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0154583647869352 lu0 = -2.91118928771256e-08 wu0 = -5.92973161822057e-09 pu0 = 2.06758831770759e-14   a0 = 1.15335206049834 la0 = -3.96226992370915e-07 wa0 = 1.06216639582676e-07 pa0 = 2.20305481552042e-14   keta = -0.033598684533428 lketa = 6.19954215161018e-08 wketa = 3.51686179093151e-08 pketa = -7.44552966088624e-14   a1 = 0.0   a2 = 0.8   ags = 0.96166140881989 lags = -2.19177842382632e-06 wags = -6.22784987229046e-07 pags = 2.08451412101801e-12   b0 = -5.5908721552003e-08 lb0 = 3.7514966807298e-13 wb0 = 4.3628493862293e-14 pb0 = -2.9274886881002e-19   b1 = -1.17955413651603e-09 lb1 = -1.10583002312134e-15 wb1 = 9.20467665449384e-16 pb1 = 8.62936891368787e-22   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.310289417538083+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.5081371230768e-07 wvoff = 7.9766557431796e-08 pvoff = -2.12747698536978e-13   nfactor = {3.36742773591543+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.34419878340445e-06 wnfactor = -8.74093743793719e-07 pnfactor = 3.19979823990222e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.16157665925 leta0 = -3.30568446409198e-7   etab = -0.141315438284516 letab = 2.8898748558036e-07 wetab = -3.46208200047724e-15 petab = 1.40291976580914e-20   dsub = 0.867836450000001 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = -2.56547909147169 lpclm = 6.29536217912578e-06 wpclm = 1.77997506938415e-06 ppclm = -3.89281872392573e-12   pdiblc1 = 0.39   pdiblc2 = 0.00567626413030715 lpdiblc2 = -1.16479175061118e-08 wpdiblc2 = -2.96065352011028e-09 ppdiblc2 = 6.41939506734754e-15   pdiblcb = 0.3705118699923 lpdiblcb = -2.41315880659321e-06 wpdiblcb = -4.64708997874606e-07 ppdiblcb = 1.88311378367438e-12   drout = 0.56   pscbe1 = 799999841.891162 lpscbe1 = 0.000324477754475083 wpscbe1 = 9.17588113225065e-05 ppscbe1 = -1.88311377775918e-10   pscbe2 = 9.65222966171759e-09 lpscbe2 = -1.50422129588033e-15 wpscbe2 = -1.18517293702406e-17 ppscbe2 = 7.49579090932929e-22   pvag = 0.0   delta = 0.01   alpha0 = -1.26270905854266e-10 lalpha0 = 2.61429922211984e-16 walpha0 = 9.60943450066332e-17 palpha0 = -1.94114130407519e-22   alpha1 = 9.9952420983626e-15 lalpha1 = -4.08985166230727e-20 walpha1 = -5.4585683026281e-21 palpha1 = 2.24279705439409e-26   beta0 = 94.9457716153883 lbeta0 = -0.000188695066177279 wbeta0 = -2.90606991709737e-05 pbeta0 = 5.96396164487366e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.10532742117647e-10 lagidl = -1.56523972879148e-15 wagidl = -5.04367041025418e-16 pagidl = 1.51640110153747e-21   bgidl = -890976974.866783 lbgidl = 3880.74425983153 wbgidl = 1475.62804248664 pbgidl = -0.00302834732079691   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.911951304157927 lkt1 = 1.02276171854909e-06 wkt1 = 3.59441477163733e-07 pkt1 = -8.2955625150524e-13   kt2 = 0.143768098117655 lkt2 = -3.17192125624822e-07 wkt2 = -1.18014499762683e-07 pkt2 = 1.86561937415698e-13   at = 156733.184894659 lat = -0.499731673046089 wat = -0.0408957945286925 pat = 2.34837141075769e-7   ute = 2.29469742402412 lute = -6.12705201394739e-06 wute = -1.18464946011941e-06 pute = 2.10415480947035e-12   ua1 = 1.35596323181477e-08 lua1 = -2.90024330500836e-14 wua1 = -7.4234708133989e-15 pua1 = 1.59059806261699e-20   ub1 = -1.19692237591462e-17 lub1 = 2.74685213997932e-23 wub1 = 7.13671316224325e-24 pub1 = -1.57172065723951e-29   uc1 = -4.81724721346144e-10 luc1 = 1.20926768082468e-15 wuc1 = 1.99889532604723e-16 puc1 = -4.83331084673622e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.85 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.819791538952487+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.62766692759225e-07 wvth0 = -1.6933153056627e-07 pvth0 = 2.15090619339543e-13   k1 = 0.635289856278905 lk1 = -2.86906578973086e-07 wk1 = -1.29561731551205e-07 pk1 = 2.11038092418321e-13   k2 = 0.00332958692698397 lk2 = -1.8191014396897e-08 wk2 = 2.80130161683075e-09 pk2 = 1.38779585377647e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 380560.359198367 lvsat = -0.545413380310392 wvsat = -0.235049432936275 pvsat = 3.84114873849229e-7   ua = -6.48738952685549e-09 lua = 8.84046946244304e-15 wua = 4.02045427203068e-15 pua = -6.40490672322082e-21   ub = 4.11213480357107e-18 lub = -4.78319468056299e-24 wub = -2.38377199780322e-24 pub = 3.53260203476338e-30   uc = 1.58334259826638e-10 luc = -2.89994835275991e-16 wuc = -1.55702628688835e-16 puc = 2.20151740193661e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.0173910136493207 lu0 = 3.83030140730315e-08 wu0 = 1.75939673112826e-08 pu0 = -2.76004632851044e-14   a0 = 2.72881387886286 la0 = -3.62945748087677e-06 wa0 = -9.45815975811675e-07 pa0 = 2.18105711886996e-12   keta = 0.150214799680107 lketa = -3.15234514766735e-07 wketa = -9.3858506016422e-08 pketa = 1.90339715277864e-13   a1 = 0.0   a2 = -0.421343079969202 la2 = 2.50649278646523e-06 wa2 = 9.53077759408742e-07 pa2 = -1.95594716020228e-12   ags = -3.22354499757013 lags = 6.39728212724275e-06 wags = 2.27468849245532e-06 pags = -3.86180554534987e-12   b0 = 4.18303565649651e-07 lb0 = -5.98049178850605e-13 wb0 = -3.2642410772255e-13 pb0 = 4.66688992424263e-19   b1 = 2.90313914113716e-08 lb1 = -6.31060315471548e-14 wb1 = -2.26547101569249e-14 pb1 = 4.92449305510917e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0769532851321222+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.28048732069527e-07 wvoff = -1.13433007816158e-07 pvoff = 1.83744756846179e-13   nfactor = {-2.62947097748348+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.96289462287749e-06 wnfactor = 2.99635800518568e-06 pnfactor = -4.74330926877852e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.16872333846843 leta0 = -2.39747816880847e-06 weta0 = -9.76904703393961e-07 peta0 = 2.00484583920733e-12   etab = -0.476090949018803 letab = 9.76028184056227e-07 wetab = 3.76465721890617e-07 petab = -7.72599135565802e-13   dsub = -0.971680209976901 ldsub = 2.52770708916362e-06 wdsub = 7.14808319556557e-07 pdsub = -1.46696037015171e-12   voffl = 0.0   minv = 0.0   pclm = 1.57613721813822 lpclm = -2.20424090095699e-06 wpclm = -9.70708286262565e-07 ppclm = 1.75225193791675e-12   pdiblc1 = 0.423414691906398 lpdiblc1 = -6.85750675620609e-08 wpdiblc1 = -1.97027859047051e-08 ppdiblc1 = 4.04349044534298e-14   pdiblc2 = 0.000431395481945641 lpdiblc2 = -8.84172536592372e-10 wpdiblc2 = -1.68864690406341e-10 ppdiblc2 = 6.89965984109438e-16   pdiblcb = -2.2371438799692 lpdiblcb = 2.93838445267503e-06 wpdiblcb = 1.40595687545358e-06 ppdiblcb = -1.95594716020228e-12   drout = 0.120527753863881 ldrout = 9.0190384082713e-07 wdrout = 5.452238580528e-08 pdrout = -1.11893184612185e-13   pscbe1 = 796324642.803025 lpscbe1 = 7.54272607998973 wpscbe1 = 2.86807307444451 ppscbe1 = -5.88598289051698e-6   pscbe2 = 1.12802684722218e-08 lpscbe2 = -4.84535254846595e-15 wpscbe2 = -6.98873784696105e-16 ppscbe2 = 2.15951529482107e-21   pvag = 0.0   delta = 0.01   alpha0 = -1.02932960431092e-10 lalpha0 = 2.13534787082894e-16 walpha0 = 3.09481647192854e-18 palpha0 = -3.25649896887149e-24   alpha1 = -1.05244685850994e-10 lalpha1 = 2.15967283973907e-16 walpha1 = 1.1225661954828e-20 palpha1 = -1.18121242123434e-26   beta0 = -6.19084066646315 lbeta0 = 1.88618384218643e-05 wbeta0 = 2.32664127452719e-06 pbeta0 = -4.7748332691595e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.40596726191037e-09 lagidl = -2.99244035399446e-15 wagidl = -7.81484020530863e-16 pagidl = 2.08511248290866e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.322737309238521 lkt1 = -1.86448578026296e-07 wkt1 = -8.04667598079586e-08 pkt1 = 7.32423484622554e-14   kt2 = 0.0577552405506807 lkt2 = -1.40672840773002e-07 wkt2 = -6.5533477591638e-08 pkt2 = 7.8858127032327e-14   at = -50008.0010014743 lat = -0.0754485214790495 wat = 0.0321252792182427 pat = 8.49801536261379e-8   ute = 2.93128622972457 lute = -7.4334869343245e-06 wute = -2.74088283575646e-06 pute = 5.29792386098787e-12   ua1 = 2.87562976713318e-09 lua1 = -7.076263602782e-15 wua1 = -2.29207719542827e-15 pua1 = 5.37511399344497e-21   ub1 = -5.51262035246808e-19 lub1 = 4.03608937765286e-24 wub1 = 1.23191012658945e-24 pub1 = -3.59911587609586e-30   uc1 = 1.79686902920536e-11 luc1 = 1.83775374644066e-16 wuc1 = 4.61036528594544e-17 puc1 = -1.67725089467553e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.86 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.20625123757844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.43882819902042e-07 wvth0 = 1.17609791292017e-07 pvth0 = -8.68413779965854e-14   k1 = 0.289168826506188 lk1 = 7.72968517580473e-08 wk1 = 8.04843601655936e-08 pk1 = -9.98143726803879e-15   k2 = -0.0378923198787193 lk2 = 2.51844484860566e-08 wk2 = 4.67871135047188e-08 pk2 = -3.24058041205823e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -355170.73772815 lvsat = 0.228754516312857 wvsat = 0.266736792513204 pvsat = -1.43886169376407e-7   ua = 3.15342462526988e-09 lua = -1.30400974343182e-15 wua = -2.69604134958043e-15 pua = 6.62478779150114e-22   ub = -8.79218610529931e-19 lub = 4.68922009950892e-25 wub = 1.08288176254463e-24 pub = -1.15160117986318e-31   uc = -1.9479040434383e-10 luc = 8.15781207247353e-17 wuc = 9.08478380285191e-17 puc = -3.92792625564077e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0253612384756981 lu0 = -6.68274395975466e-09 wu0 = -1.24024013446698e-08 pu0 = 3.96300565854084e-15   a0 = -2.86976139471617 la0 = 2.26160416071985e-06 wa0 = 2.44943864711099e-06 pa0 = -1.39157579131806e-12   keta = -0.200071965391825 lketa = 5.33522817728494e-08 wketa = 1.22732770790608e-07 pketa = -3.75669396033951e-14   a1 = 0.0   a2 = 3.2426861599384 la2 = -1.34895633302286e-06 wa2 = -1.90615551881748e-06 pa2 = 1.05266104217832e-12   ags = 3.02515908547085 lags = -1.77873003208538e-07 wags = -1.73818977105249e-06 pags = 3.60717517278382e-13   b0 = -5.40461278333841e-07 lb0 = 4.10804416877117e-13 wb0 = 4.21750147562625e-13 pb0 = -3.20572130479776e-19   b1 = -6.56683122489154e-08 lb1 = 3.65410687314565e-14 wb1 = 5.12444119337281e-14 pb1 = -2.85149033749433e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.371530090376825+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 8.19176492115754e-08 wvoff = 1.14667010569041e-07 pvoff = -5.62718907995182e-14   nfactor = {5.98933445540839+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.10618306224496e-06 wnfactor = -2.98520287742129e-06 pnfactor = 1.5507462990185e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -2.87659257393686 leta0 = 1.85917718280861e-06 weta0 = 1.95380940678792e-06 peta0 = -1.07897756823278e-12   etab = 0.950136534213168 letab = -5.24709701582233e-07 wetab = -7.52931429932906e-07 petab = 4.15801111660438e-13   dsub = 2.59657816045177 ldsub = -1.22696780331135e-06 wdsub = -1.38017012747168e-06 pdsub = 7.37466035884625e-13   voffl = 0.0   minv = 0.0   pclm = -1.76881329444398 lpclm = 1.31545986125403e-06 wpclm = 1.45044922444083e-06 ppclm = -7.95394104618328e-13   pdiblc1 = 0.714029335749044 lpdiblc1 = -3.74372292242979e-07 wpdiblc1 = -6.3188896424419e-08 ppdiblc1 = 8.61928598450252e-14   pdiblc2 = -0.000152581521148273 lpdiblc2 = -2.69686822925823e-10 wpdiblc2 = 1.34588293737908e-11 ppdiblc2 = 4.98117336685433e-16   pdiblcb = 0.5553522 wpdiblcb = -4.5287911604484e-7   drout = 0.425392371916349 ldrout = 5.81112180533744e-07 wdrout = 3.02652100137375e-07 pdrout = -3.72985939610132e-13   pscbe1 = 807350714.393948 lpscbe1 = -4.05938056905734 wpscbe1 = -5.73614614888947 ppscbe1 = 3.16774655770118e-6   pscbe2 = -2.28982905519193e-08 lpscbe2 = 3.11187969347734e-14 wpscbe2 = 2.36493987282457e-14 ppscbe2 = -2.34607840190144e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 14.8063323637092 lbeta0 = -3.23228991892331e-06 wbeta0 = -4.72100369308145e-06 pbeta0 = 2.64100181449191e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -3.60392094320944e-09 lagidl = 2.27917944062543e-15 wagidl = 2.65044333818453e-15 pagidl = -1.5261090568081e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.493519010598582 lkt1 = -6.74472824207854e-09 wkt1 = -2.05055389328904e-08 pkt1 = 1.01485735250111e-14   kt2 = -0.164265742222121 lkt2 = 9.2947184202799e-08 wkt2 = 7.08522414834577e-08 pkt2 = -6.4652791164409e-14   at = -325045.311993826 lat = 0.213957563751476 wat = 0.235316613718021 pat = -1.28826505761912e-7   ute = -7.95606229665975 lute = 4.02264934112371e-06 wute = 4.45602556453441e-06 pute = -2.2749726248594e-12   ua1 = -9.49643456110342e-09 lua1 = 5.94215448215466e-15 wua1 = 6.53627574458814e-15 pua1 = -3.91445858921672e-21   ub1 = 6.06405519451678e-18 lub1 = -2.92483187014527e-24 wub1 = -4.41929511307645e-24 pub1 = 2.3473252789059e-30   uc1 = 3.78504506926095e-10 luc1 = -1.95595914658387e-16 wuc1 = -2.38425686943524e-16 puc1 = 1.31668916634753e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.87 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.897664768814751+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.65318973674235e-08 wvth0 = -8.75687760964322e-08 pvth0 = 2.64670495937139e-14   k1 = 0.246452479905976 lk1 = 1.00886655153588e-07 wk1 = 1.37861948971556e-07 pk1 = -4.166780904301e-14   k2 = 0.0474129623487683 lk2 = -2.19247964870978e-08 wk2 = -2.62717927895834e-08 pk2 = 7.94046546810206e-15   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 23344.8119907215 lvsat = 0.0197219535894583 wvsat = 0.0136694285258487 pvsat = -4.13148908593808e-9   ua = 3.55690043806238e-09 lua = -1.52682643671579e-15 wua = -3.30556473546492e-15 pua = 9.99083802341123e-22   ub = -1.75679650814316e-18 lub = 9.53558260862512e-25 wub = 1.93141502082646e-24 pub = -5.83756670139652e-31   uc = -1.04041082279571e-10 luc = 3.14624428600023e-17 wuc = 4.35632802399032e-17 puc = -1.31666965095491e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0237376109832811 lu0 = -5.78610704245984e-09 wu0 = -1.15445346689745e-08 pu0 = 3.48925479195486e-15   a0 = 1.72537582435042 la0 = -2.76028202549144e-07 wa0 = -1.55561778086173e-07 pa0 = 4.70174584940991e-14   keta = -0.21649122006379 lketa = 6.24197002306592e-08 wketa = 1.2084549574529e-07 pketa = -3.65247051705436e-14   a1 = 0.0   a2 = 1.13401084291128 la2 = -1.84455149921854e-7   ags = 5.46105100897625 lags = -1.52307726672093e-06 wags = -2.39674246582784e-06 pags = 7.24398633099204e-13   b0 = 4.49353836584809e-07 lb0 = -1.35814051630902e-13 wb0 = -3.50654254957396e-13 pb0 = 1.05982793981088e-19   b1 = 1.10481188071491e-09 lb1 = -3.33921657262918e-16 wb1 = -8.62142381702021e-16 pb1 = 2.60576499872764e-22   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.251959941063855+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.58858712445328e-08 wvoff = 2.82086524726427e-08 pvoff = -8.52586774928903e-15   nfactor = {2.08960844309255+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 4.74133299743794e-08 wnfactor = -3.91244374469089e-07 pnfactor = 1.18250873472661e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.1754675e-05 letab = -3.7555105736025e-11 wetab = 1.29246970711411e-26 petab = 3.08148791101958e-33   dsub = 0.0686624724021905 ldsub = 1.69055940004215e-07 wdsub = -9.88930232828686e-08 pdsub = 2.98897240360841e-14   voffl = 0.0   minv = 0.0   pclm = 0.584279929133476 lpclm = 1.59806001859505e-08 wpclm = 2.24253057382051e-08 ppclm = -6.77789168223234e-15   pdiblc1 = -0.478703349304998 lpdiblc1 = 2.8430598394932e-07 wpdiblc1 = 2.05188936467658e-07 ppdiblc1 = -6.20169197247945e-14   pdiblc2 = -0.0147960134174852 lpdiblc2 = 7.81704593780299e-09 wpdiblc2 = 2.02219952398121e-09 ppdiblc2 = -6.11195650726654e-16   pdiblcb = 1.4987761599384 lpdiblcb = -5.20999277908262e-07 wpdiblcb = -1.0003972867278e-06 ppdiblcb = 3.02363077132471e-13   drout = 2.7422400234303 ldrout = -6.98350717081274e-07 wdrout = -8.23393743495871e-07 pdrout = 2.48864995215423e-13   pscbe1 = 800086006.26808 lpscbe1 = -0.0474963595029294   pscbe2 = 6.27592696057523e-08 lpscbe2 = -1.61849910593797e-14 wpscbe2 = -4.16022764685272e-14 ppscbe2 = 1.25739968466771e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.54244020089537 lbeta0 = 2.26900680745475e-07 wbeta0 = 1.35442288054147e-07 pbeta0 = -4.09364834683496e-14   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.03486010873846e-09 lagidl = -2.82554923845438e-16 wagidl = -2.49681105596234e-16 pagidl = 7.54643663987225e-23   bgidl = 664683394.790398 lbgidl = 185.176248010765   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.49807029680829 lkt1 = -4.23131229177233e-09 wkt1 = -4.70186724762058e-09 pkt1 = 1.42110646252255e-15   kt2 = 0.0301985471073132 lkt2 = -1.44443583293557e-08 wkt2 = -1.0210054708344e-07 pkt2 = 3.085917565214e-14   at = 57349.9216482771 lat = 0.00278247273925974 wat = 0.0045017877902751 pat = -1.36063384709613e-9   ute = -1.26013523664223 lute = 3.24870493718457e-07 wute = 7.43345203903094e-07 pute = -2.24670884463283e-13   ua1 = 2.30460029442892e-09 lua1 = -5.74884409569079e-16 wua1 = -1.21938425279252e-15 pua1 = 3.68550354716769e-22   ub1 = 1.16526194256105e-18 lub1 = -2.19507588305478e-25 wub1 = -3.72798048899116e-25 pub1 = 1.12675600693416e-31   uc1 = 5.303025600552e-11 luc1 = -1.58550379072564e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.88 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.25148808693957+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 8.04087237725772e-08 wvth0 = 2.03910099959358e-07 pvth0 = -6.1630400342016e-14   k1 = -2.64769270144974 lk1 = 9.75621777202084e-07 wk1 = 1.09909331904171e-06 pk1 = -3.32193262027124e-13   k2 = 0.994001379408727 lk2 = -3.08024519424551e-07 wk2 = -2.63285938358031e-07 pk2 = 7.95763318671464e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -40614.912625554 lvsat = 0.0390533326366552 wvsat = 0.0157316243944771 pvsat = -4.75477335185991e-9   ua = 1.2051495474672e-09 lua = -8.16026192289627e-16 wua = 2.47015051308807e-16 pua = -7.46585701527286e-23   ub = -1.62828057149119e-18 lub = 9.14715218621011e-25 wub = 4.11055926101477e-25 pub = -1.24238776272689e-31   uc = -2.0014119224054e-12 luc = 6.21666772241634e-19 wuc = 1.15533172761559e-18 puc = -3.49190927349718e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00785199502177666 lu0 = -9.84790817406843e-10 wu0 = 2.51794640344037e-09 pu0 = -7.61031674815027e-16   a0 = 1.95745393042207 la0 = -3.46172185562559e-07 wa0 = -1.60546711227303e-06 pa0 = 4.85241196414739e-13   keta = 0.187099559975319 lketa = -5.95627879007013e-08 wketa = -2.49816505023507e-07 pketa = 7.550528992782e-14   a1 = 0.0   a2 = -0.192308203327515 la2 = 2.16415497570498e-07 wa2 = 1.36582654162594e-07 pa2 = -4.12811511420647e-14   ags = -2.32595109449885 lags = 8.30489610039698e-7   b0 = -6.79767101600045e-07 lb0 = 2.05454848088903e-13 wb0 = 5.30457753221219e-13 pb0 = -1.60327142706841e-19   b1 = 3.3314441400079e-09 lb1 = -1.00690567120841e-15 wb1 = -2.59969976383228e-15 pb1 = 7.85741055719959e-22   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.339380792821851+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.62842726187285e-07 wvoff = -3.07029470449379e-07 pvoff = 9.27975082370315e-14   nfactor = {-1.3206882242339+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.07815162559713e-06 wnfactor = 3.80462724791569e-06 pnfactor = -1.14992195329178e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.570090261060969 leta0 = -2.42067207738505e-08 weta0 = 6.58881148553885e-07 peta0 = -1.99142214982372e-13   etab = -0.543821641413894 letab = 1.6434739417836e-07 wetab = 5.05857714813868e-07 petab = -1.52891953298488e-13   dsub = 1.73672279469971 ldsub = -3.35103615987956e-07 wdsub = 6.3002901885497e-08 pdsub = -1.90421860745781e-14   voffl = 0.0   minv = 0.0   pclm = 0.725036330252816 lpclm = -2.65620367575624e-08 wpclm = -2.95003267155116e-08 ppclm = 8.91626724747629e-15   pdiblc1 = 1.65229349989834 lpdiblc1 = -3.59772896744446e-07 wpdiblc1 = -1.270473665246e-07 ppdiblc1 = 3.83991772004948e-14   pdiblc2 = 0.0503771960865463 lpdiblc2 = -1.1881100422324e-08 wpdiblc2 = -8.01493282081463e-09 ppdiblc2 = 2.42245734056148e-15   pdiblcb = -0.000668890291118274 lpdiblcb = -6.78025075917416e-08 wpdiblcb = -5.6341013781391e-07 ppdiblcb = 1.70286770283289e-13   drout = -1.453869509709 ldrout = 5.69894016543347e-7   pscbe1 = 799692834.756853 lpscbe1 = 0.0713369775635329   pscbe2 = -7.21404676956558e-08 lpscbe2 = 2.45875102418098e-14 wpscbe2 = 6.30191902020444e-14 ppscbe2 = -1.90471091042365e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.94818744040796 lbeta0 = 7.08752417833477e-07 wbeta0 = 3.12646576909388e-06 pbeta0 = -9.44952393448243e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.35724510864813e-08 lagidl = -1.31392440337314e-14 wagidl = -3.3923822844728e-14 pagidl = 1.02532379880591e-20   bgidl = 2159327259.4845 lbgidl = -266.569397585975 wbgidl = 22.1880513307788 pbgidl = -6.70618319836835e-6   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.055031774217257 lkt1 = -1.71402541544746e-07 wkt1 = -1.16296822171205e-07 pkt1 = 3.51499004234915e-14   kt2 = 0.322172873485714 lkt2 = -1.02691554656943e-07 wkt2 = -2.64697796016969e-23 pkt2 = -6.31088724176809e-30   at = 438135.742396925 lat = -0.112307376081274 wat = -0.27077325999319 pat = 8.18393224201218e-8   ute = 0.726393300964688 lute = -2.7554385107347e-07 wute = -6.31443663016137e-07 pute = 1.90849427040987e-13   ua1 = 1.38344640470347e-09 lua1 = -2.9647209447679e-16 wua1 = -1.12916100596461e-16 pua1 = 3.41281009925762e-23   ub1 = -1.99870168567005e-19 lub1 = 1.93094036358197e-25 wub1 = 4.98543741555632e-25 pub1 = -1.50681356078999e-31   uc1 = 2.24422226624312e-10 luc1 = -6.7657061282992e-17 wuc1 = -1.75637125429771e-16 puc1 = 5.30850917012702e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.89 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.0931089549404156+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.31864527024756e-07 wvth0 = -7.05288330146851e-07 pvth0 = 1.4952457066114e-13   k1 = 2.80462855665424 lk1 = -2.90641668743759e-07 wk1 = -2.42375184290739e-06 pk1 = 4.85962866919423e-13   k2 = -0.370820399272816 lk2 = 8.94578492178751e-09 wk2 = 5.44429902117225e-07 pk2 = -1.08010018072348e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1169817.44248675 lvsat = -0.242061108811692 wvsat = -0.46580046642803 pvsat = 1.07077684017032e-7   ua = 7.70293651976377e-10 lua = -7.15033954553152e-16 wua = -1.7074029745474e-15 pua = 3.79241335426195e-22   ub = -2.50706242416423e-18 lub = 1.11880615243135e-24 wub = 2.63723016485163e-24 pub = -6.4125216000274e-31   uc = 3.97535127112923e-12 luc = -7.6639464211443e-19 wuc = -2.53025421502165e-18 puc = 5.06760608726183e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00597068720161809 lu0 = -5.47870245329753e-10 wu0 = -1.53162782409541e-09 pu0 = 1.79453592510567e-16   a0 = -3.23502716693098 la0 = 8.59745201930004e-07 wa0 = 3.58174859154209e-06 pa0 = -7.19453340286396e-13   keta = -3.08184186925686 lketa = 6.99625976448467e-07 wketa = 2.06041001348967e-06 pketa = -4.61028647411235e-13   a1 = 0.0   a2 = -1.01295383316313 la2 = 4.07004700580411e-07 wa2 = -3.18692859712718e-07 pa2 = 6.44534000268795e-14   ags = 18.9018185895908 lags = -4.09951130470234e-06 wags = -1.02442717524699e-05 pags = 2.37916040460888e-12   b0 = 2.71545869463027e-06 lb0 = -5.83062576505014e-13 wb0 = -2.11901416636386e-12 pb0 = 4.54994164313356e-19   b1 = 2.81059978643752e-07 lb1 = -6.55074137099614e-14 wb1 = -2.19325772666605e-13 pb1 = 5.11188544048785e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.97195323274911+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 6.06191421913393e-07 wvoff = 2.39345982250479e-06 pvoff = -5.34372226626522e-13   nfactor = {13.9587862778434+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -2.47039937118881e-06 wnfactor = -5.62061783047231e-06 pnfactor = 1.03902523944828e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.145259210231043 leta0 = 1.4192818648742e-07 weta0 = -7.22355569432068e-07 peta0 = 1.2164034411284e-13   etab = 2.36021930674408 letab = -5.10095787744692e-07 wetab = -1.81403969977418e-06 petab = 3.85887981957684e-13   dsub = 0.615654716810817 ldsub = -7.47434023748049e-08 wdsub = -2.2022267849703e-07 pdsub = 4.67349723902009e-14   voffl = 0.0   minv = 0.0   pclm = 1.57856979309032 lpclm = -2.24789208767333e-07 wpclm = 1.02499210535736e-06 ppclm = -2.35982218654425e-13   pdiblc1 = 0.47650235885655 lpdiblc1 = -8.67036347754758e-08 wpdiblc1 = 4.45280255706734e-07 ppdiblc1 = -9.45199067693772e-14   pdiblc2 = -0.0131496281443229 lpdiblc2 = 2.87255981752574e-09 wpdiblc2 = 2.1983543361775e-08 ppdiblc2 = -4.54447876351169e-15   pdiblcb = -2.38502081431666 lpdiblcb = 4.85946536299721e-07 wpdiblcb = 1.40820633441033e-06 ppdiblcb = -2.87607354075485e-13   drout = 1.0   pscbe1 = 1613549587.36535 lpscbe1 = -188.941196818491 wpscbe1 = -472.017318047236 ppscbe1 = 0.000109622717995244   pscbe2 = 2.06347087681145e-07 lpscbe2 = -4.00892750815645e-14 wpscbe2 = -1.50609837883802e-13 ppscbe2 = 3.05667372655048e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 37.2499460182054 lbeta0 = -6.32861889954995e-06 wbeta0 = -1.4149754088154e-05 pbeta0 = 3.06732873485857e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -7.27680961892001e-08 lagidl = 1.38800336872147e-14 wagidl = 5.62242639543309e-14 pagidl = -1.06830241344147e-20   bgidl = 1089208104.61615 lbgidl = -18.0417147018843 wbgidl = -51.7721197718129 pbgidl = 1.04705488190109e-5   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.502593517506934 lkt1 = -4.18979709188448e-08 wkt1 = 2.71359251732812e-07 pkt1 = -5.48805091481993e-14   kt2 = -0.12   at = -89229.7398926124 lat = 0.0101695656220953 wat = 0.315874207226237 pat = -5.44054453093195e-8   ute = -1.5255072250135 lute = 2.47444282781283e-07 wute = 1.00212960520176e-06 pute = -1.88536529489744e-13   ua1 = 1.41338028698651e-09 lua1 = -3.03424029099851e-16 wua1 = -7.59912923055232e-16 pua1 = 1.84388584030868e-22   ub1 = 2.40220412232301e-18 lub1 = -4.11219503180973e-25 wub1 = -1.16326873029648e-24 pub1 = 2.3526295782135e-31   uc1 = -5.71554220936062e-10 luc1 = 1.17202896827772e-16 wuc1 = 4.09819959336132e-16 puc1 = -8.28832180360174e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.90 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0283044+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47866595   k2 = 0.0129645355   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24491.02   ua = -9.0471719e-10   ub = 6.9558965e-19   uc = -6.8009552e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0063669233   a0 = 1.2509318   keta = 0.0074076058   a1 = 0.0   a2 = 0.8   ags = 0.23496304   b0 = 3.1294e-9   b1 = 2.2449e-9   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20719556+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4509367+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00083787503   pdiblcb = -0.225   drout = 0.56   pscbe1 = 790097310.0   pscbe2 = 9.5178184e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1731672e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.52561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.91 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0283044+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47866595   k2 = 0.0129645355   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24491.02   ua = -9.0471719e-10   ub = 6.9558965e-19   uc = -6.8009552e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0063669233   a0 = 1.2509318   keta = 0.0074076058   a1 = 0.0   a2 = 0.8   ags = 0.23496304   b0 = 3.1294e-9   b1 = 2.2449e-9   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20719556+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4509367+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00083787503   pdiblcb = -0.225   drout = 0.56   pscbe1 = 790097310.0   pscbe2 = 9.5178184e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1731672e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.52561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.92 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.03539511610748+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.70961691413993e-8   k1 = 0.495157110071913 lk1 = -1.32790828250936e-7   k2 = 0.00836364767003139 lk2 = 3.70474668226501e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -7382.89011603501 lvsat = 0.256656469614472   ua = -9.58466181674431e-10 lua = 4.32799941967484e-16   ub = 7.6909750010972e-19 lub = -5.91903071491038e-25   uc = -6.32758098636854e-11 luc = -3.81172419809453e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00587902240304999 lu0 = 3.92869658215954e-9   a0 = 1.25394119826395 la0 = -2.42324061051148e-8   keta = 0.0041337224981316 lketa = 2.63621039002867e-8   a1 = 0.0   a2 = 0.8   ags = 0.235897132664538 lags = -7.52154111937366e-9   b0 = 1.91017210088e-08 lb0 = -1.28613010036863e-13 wb0 = 3.15544362088405e-30 pb0 = -1.20370621524202e-35   b1 = 4.01204264987e-09 lb1 = -1.42294620324172e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.213052925297388+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.71649287143317e-8   nfactor = {0.992893134698274+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.68827809239585e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.40154855792662 lpclm = 3.24737935499048e-06 wpclm = 4.79764755280756e-23 ppclm = -2.08259278978347e-28   pdiblc1 = 0.39   pdiblc2 = 0.00125107721379807 lpdiblc2 = -3.32720439207274e-09 wpdiblc2 = -8.27180612553028e-25   pdiblcb = -0.225   drout = 0.56   pscbe1 = 780065283.441584 lpscbe1 = 80.7803156308364   pscbe2 = 9.4554969287815e-09 lpscbe2 = 5.01827630368908e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.79745850696584e-10 lalpha0 = -6.4213296805061e-16   alpha1 = 2.0130604093734e-10 lalpha1 = -8.15740858995407e-16   beta0 = -17.9357625134483 lbeta0 = 0.000168579847148576 pbeta0 = -2.58493941422821e-26   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.2603507685074e-09 lagidl = -8.75426627922873e-15   bgidl = 674167346.162077 lbgidl = 2623.68370603786   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.660002639095 lkt1 = 1.08216218740424e-6   kt2 = -0.0463613991892905 lkt2 = -4.93006695198299e-8   at = -43490.6338305398 lat = 0.430719581827527 pat = 5.29395592033938e-23   ute = -2.1668478607375 lute = 7.3061854601885e-6   ua1 = -8.95048198670001e-10 lua1 = 5.14536877225312e-15   ub1 = 5.6628226602667e-19 lub1 = -5.79296608017391e-25   uc1 = 6.14761923450098e-11 luc1 = -4.29032302867458e-16 wuc1 = -6.16297582203915e-33 puc1 = 4.70197740328915e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.93 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.982614265333149+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.56784663942897e-7   k1 = 0.47568105030166 lk1 = -5.38691013793489e-8   k2 = 0.024238964229633 lk2 = -2.72831735787798e-08 wk2 = 1.32348898008484e-23   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 80233.7862794006 lvsat = -0.0983875939921968   ua = -1.07940391206423e-09 lua = 9.22869013375441e-16   ub = 6.05632862096945e-19 lub = 7.04953636437602e-26   uc = -7.91086515473494e-11 luc = 2.60412799017912e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00524089405412752 lu0 = 6.51454771718224e-9   a0 = 1.3363730597858 la0 = -3.58266339933986e-7   keta = 0.0270000655175154 lketa = -6.62978745356101e-8   a1 = 0.0   a2 = 0.8   ags = -0.111454170356075 lags = 1.40003034508678e-06 pags = 4.03896783473158e-28   b0 = 1.9267169678e-08 lb0 = -1.29283448248488e-13 pb0 = -2.40741243048404e-35   b1 = 4.06495964525e-10 lb1 = 3.81089284445321e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17284433258485+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.15770059644899e-7   nfactor = {1.8612841496695+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.69346680715817e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.16157665925 leta0 = -3.30568446409198e-7   etab = -0.14131544425 letab = 2.88987509753953e-7   dsub = 0.86783645 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = 0.50158099615122 lpclm = -4.12321058614568e-7   pdiblc1 = 0.39   pdiblc2 = 0.000574786923689725 lpdiblc2 = -5.86711798013223e-10   pdiblcb = -0.4302243 lpdiblcb = 8.31618733104899e-7   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.63180804641184e-09 lpscbe2 = -2.12627861870897e-16   pvag = 0.0   delta = 0.01   alpha0 = 3.93084526915155e-11 lalpha0 = -7.30465050463587e-17   alpha1 = 5.89628916180988e-16 lalpha1 = -2.25306900705458e-21 walpha1 = -9.4039548065783e-38 palpha1 = 2.69049305150365e-43   beta0 = 44.8715250268964 lbeta0 = -8.59305441357732e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.58537868841385e-10 lagidl = 1.04765826924742e-15 pagidl = 1.88079096131566e-37   bgidl = 1651665307.67585 lbgidl = -1337.37556602061   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.292600714699091 lkt1 = -4.06639688915615e-7   kt2 = -0.0595816949264356 lkt2 = 4.27118133894581e-9   at = 86265.9849276524 lat = -0.0950857682390263 wat = -5.55111512312578e-17   ute = 0.253437892106421 lute = -2.501400539773e-06 pute = -8.07793566946316e-28   ua1 = 7.68312127754843e-10 lua1 = -1.59497146697967e-15   ub1 = 3.2798673173032e-19 lub1 = 3.86334802766253e-25   uc1 = -1.37296747083752e-10 luc1 = 3.76443949522164e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.94 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.111565276635+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.07854146344242e-7   k1 = 0.412043125153901 lk1 = 7.6731385039666e-8   k2 = 0.008156486207853 lk2 = 5.72197936407216e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -24451.343929966 lvsat = 0.116451731684064   ua = 4.40221451496412e-10 lua = -2.19577150161434e-15 pua = 7.52316384526264e-37   ub = 4.67730137977917e-21 lub = 1.30380220643664e-24   uc = -1.09955631533875e-10 luc = 8.93467786502783e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.012925003609307 lu0 = -9.25511232866804e-9   a0 = 1.0990863172 la0 = 1.28703716530523e-7   keta = -0.0115120034860086 lketa = 1.27382494923889e-8   a1 = 0.0   a2 = 1.2208972 la2 = -8.637833324196e-7   ags = 0.69595163301957 lags = -2.56962563050263e-07 wags = -4.2351647362715e-22   b0 = -1.4415507192e-07 lb0 = 2.06098703115317e-13 pb0 = -4.81482486096809e-35   b1 = -1.000474932683e-08 lb1 = 2.17474945549116e-14 wb1 = -2.36658271566304e-30 pb1 = -3.76158192263132e-36   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.27240874789449+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 8.85603147234018e-8   nfactor = {2.5335283273967+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.21026172731559e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.5145729485 leta0 = 1.05705485304849e-06 weta0 = -3.35008148083976e-23 peta0 = 1.69605094622518e-28   etab = 0.1725939735 letab = -3.55230895457561e-07 wetab = 3.35008148083976e-23 petab = 3.23432971140615e-29   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = -0.09648207453021 lpclm = 8.15049691749903e-7   pdiblc1 = 0.38946498704665 lpdiblc1 = 1.09797658842124e-9   pdiblc2 = 0.00014042615262055 lpdiblc2 = 3.04702053888095e-10   pdiblcb = 0.1854486 lpdiblcb = -4.318916662098e-7   drout = 0.21447481877598 ldrout = 7.09101634490726e-7   pscbe1 = 801266595.421528 lpscbe1 = -2.59936158766686   pscbe2 = 1.00760449253892e-08 lpscbe2 = -1.124309887094e-15   pvag = 0.0   delta = 0.01   alpha0 = -9.7600308169365e-11 lalpha0 = 2.07923541069057e-16 walpha0 = -1.84889274661175e-32 palpha0 = 1.46936793852786e-38   alpha1 = -1.05225343007191e-10 lalpha1 = 2.15946930601916e-16 walpha1 = 1.61164977475139e-32 palpha1 = -8.63684142773358e-39   beta0 = -2.1818246335659 lbeta0 = 1.06343633314632e-05 pbeta0 = -3.23117426778526e-27   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.93987117595102e-11 lagidl = 6.00399447265296e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.46138890702338 lkt1 = -6.02453027354373e-8   kt2 = -0.055164944108976 lkt2 = -4.79306460892984e-9   at = 5346.79771944496 lat = 0.0709800672747071   ute = -1.79150595708278 lute = 1.6953211601186e-6   ua1 = -1.07382919145829e-09 lua1 = 2.18555016038624e-15 wua1 = 7.39557098644699e-32 pua1 = -7.05296610493373e-38   ub1 = 1.57143195400566e-18 lub1 = -2.16551695053176e-24 pub1 = -7.00649232162409e-46   uc1 = 9.74095071950557e-11 luc1 = -1.05230317877739e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.95 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0035987943+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.75282892738461e-9   k1 = 0.427850751319419 lk1 = 6.00979210603795e-8   k2 = 0.0427261623200538 lk2 = -3.06537203372584e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 104441.18846633 lvsat = -0.0191745332822115   ua = -1.4921015734426e-09 lua = -1.62498124883438e-16   ub = 9.86685856696402e-19 lub = 2.7049057816461e-25   uc = -3.825125789359e-11 luc = 1.38963534179038e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00399076491728 lu0 = 1.45877795346538e-10   a0 = 1.3508457592 la0 = -1.36208393997886e-7   keta = 0.0114078408200021 lketa = -1.13789962397007e-08 wketa = 8.27180612553028e-25 pketa = -1.57772181044202e-30   a1 = 0.0   a2 = -0.0417944000000006 la2 = 4.648750648392e-7   ags = 0.0300988943446807 lags = 4.4367632025122e-7   b0 = 1.86252857604e-07 lb0 = -1.41570727870806e-13   b1 = 2.263050342496e-08 lb1 = -1.25927217063902e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17394832783842+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.50439730576573e-8   nfactor = {0.845556457459399+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.65894857022848e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -0.3472332869625 letab = 1.91753700573282e-7   dsub = 0.218418609283221 ldsub = 4.37537273119964e-8   voffl = 0.0   minv = 0.0   pclm = 0.730443578263381 lpclm = -5.50770379225833e-8   pdiblc1 = 0.605149079200659 lpdiblc1 = -2.2585409959199e-07 wpdiblc1 = -4.2351647362715e-22   pdiblc2 = -0.00012939072532844 lpdiblc2 = 5.88614974991774e-10 ppdiblc2 = 1.97215226305253e-31   pdiblcb = -0.225   drout = 0.94688966293614 ldrout = -6.15767583728937e-8   pscbe1 = 797466809.156939 lpscbe1 = 1.39893691074485   pscbe2 = 1.78517897066646e-08 lpscbe2 = -9.30628290297759e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.6716105635998 lbeta0 = 1.31839811929197e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 9.63035705157761e-10 lagidl = -3.50446253579057e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.52885193245688 lkt1 = 1.07421935357837e-8   kt2 = -0.0421808401859821 lkt2 = -1.84554970731727e-8   at = 80426.768094818 lat = -0.00802230599298659   ute = -0.277922083640114 lute = 1.02663124375668e-7   ua1 = 1.7661672599772e-09 lua1 = -8.02816225661589e-16   ub1 = -1.55079508618596e-18 lub1 = 1.11982459692059e-24 pub1 = -3.50324616081204e-46   uc1 = -3.23247911165834e-11 luc1 = 3.12816893805954e-17 wuc1 = -3.08148791101958e-33   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.96 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0485537911988+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.90732534249986e-8   k1 = 0.484001245933841 lk1 = 2.90892034630282e-8   k2 = 0.0021442569150964 lk2 = -8.2426471507085e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 46898.4894401199 lvsat = 0.0126030194561198   ua = -2.1388903859664e-09 lua = 1.94686469311144e-16   ub = 1.5712084874896e-18 lub = -5.23079530325195e-26   uc = -2.89775600944163e-11 luc = 8.77501872419472e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00384532028640001 lu0 = 2.26198574637605e-10   a0 = 1.45732863148 la0 = -1.9501281483441e-7   keta = -0.00826336162663802 lketa = -5.15712386960851e-10   a1 = 0.0   a2 = 1.13401084291128 la2 = -1.84455149921854e-7   ags = 1.33124420230292 lags = -2.74872068051562e-07 wags = 8.470329472543e-22   b0 = -1.54855564116e-07 lb0 = 4.68040102651122e-14   b1 = -3.8073841392e-10 lb1 = 1.15075520438423e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.2033538489828+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.19502015567843e-9   nfactor = {1.4154585484784+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.51170416572243e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.1754675e-05 letab = -3.7555105736025e-11 petab = -1.07852076885685e-32   dsub = -0.10173926516832 ldsub = 2.20558672372739e-7   voffl = 0.0   minv = 0.0   pclm = 0.622920785045119 lpclm = 4.30167197264786e-9   pdiblc1 = -0.12514401676924 lpdiblc1 = 1.77445150605715e-7   pdiblc2 = -0.0113115784071911 lpdiblc2 = 6.76389984698667e-09 wpdiblc2 = -1.65436122510606e-24 ppdiblc2 = -3.94430452610506e-31   pdiblcb = -0.225   drout = 1.32345718174232 ldrout = -2.69533534660974e-07 wdrout = 8.470329472543e-22   pscbe1 = 800086006.268082 lpscbe1 = -0.0474963595033842   pscbe2 = -8.9252634562868e-09 lpscbe2 = 5.48115726689019e-15 wpscbe2 = -7.88860905221012e-31   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.77581966952519 lbeta0 = 1.56363370008396e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.0463669337752e-10 lagidl = -1.52522908116502e-16 pagidl = -9.4039548065783e-38   bgidl = 664683394.790401 lbgidl = 185.176248010765   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.50617204476 lkt1 = -1.78261568560315e-9   kt2 = -0.145730047776 lkt2 = 3.87288279739616e-8   at = 65106.9143680001 lat = 0.000437975988672568   ute = 0.0207166389999998 lute = -6.22580197312769e-8   ua1 = 2.0348953308e-10 lua1 = 6.01616102733013e-17   ub1 = 5.2289675656e-19 lub1 = -2.53572073929646e-26   uc1 = 5.303025600552e-11 luc1 = -1.58550379072564e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.97 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.900132306847144+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.57861012698995e-8   k1 = -0.753854237424431 lk1 = 4.03222358319681e-7   k2 = 0.540335591016728 lk2 = -1.70907210543588e-07 wk2 = -5.29395592033938e-23 pk2 = -2.52435489670724e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -13507.8828004287 lvsat = 0.03086042262122   ua = 1.63077910708428e-09 lua = -9.44669747276974e-16   ub = -9.19993558705716e-19 lub = 7.00640427015691e-25   uc = -1.06695290525573e-14 luc = 1.9978819047491e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0121906473150571 lu0 = -2.29611810248482e-9   a0 = -0.808912962428572 la0 = 4.89942843233298e-7   keta = -0.243357161001197 lketa = 7.0539742817404e-08 wketa = 2.64697796016969e-23 pketa = 1.26217744835362e-29   a1 = 0.0   a2 = 0.0430362205630015 la2 = 1.45284292860557e-7   ags = -2.32595109449885 lags = 8.30489610039698e-7   b0 = 2.34260196342857e-07 lb0 = -7.08035045232541e-14   b1 = -1.14807668171428e-09 lb1 = 3.46998140511371e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.189659108206143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.94411938088092e-9   nfactor = {5.23503302213285+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.03269231068501e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.70540283255443 leta0 = -3.67346998319748e-7   etab = 0.327817537026142 letab = -9.90994460308925e-08 wetab = 1.96455395481344e-24 petab = -2.487377041775e-29   dsub = 1.84528256562071 ldsub = -3.67915046830431e-7   voffl = 0.0   minv = 0.0   pclm = 0.674204565135856 lpclm = -1.11984915733173e-8   pdiblc1 = 1.43337925002628 lpdiblc1 = -2.93607597120365e-7   pdiblc2 = 0.0365667326803342 lpdiblc2 = -7.70698453104026e-9   pdiblcb = -0.971476165276739 lpdiblcb = 2.25617195621737e-7   drout = -1.453869509709 ldrout = 5.69894016543347e-7   pscbe1 = 799692834.756855 lpscbe1 = 0.0713369775630781   pscbe2 = 3.64473694867386e-08 lpscbe2 = -8.23240343170861e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 12.33537434018 lbeta0 = -9.1948711231432e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.48814030467986e-08 lagidl = 4.52802420107354e-15 wagidl = -7.88860905221012e-31 pagidl = -1.45761299501964e-36   bgidl = 2197559304.32 lbgidl = -278.12476551319   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.145358303 lkt1 = -1.10836043436371e-7   kt2 = 0.322172873485714 lkt2 = -1.02691554656943e-07 wkt2 = 5.29395592033938e-23 pkt2 = -2.52435489670724e-29   at = -28431.3869999999 lat = 0.028709272809041   ute = -0.361641969714285 lute = 5.33071932423549e-8   ua1 = 1.18888162042857e-09 lua1 = -2.37666250383193e-16   ub1 = 6.59166363999998e-19 lub1 = -6.65437423544523e-26   uc1 = -7.82166285911428e-11 luc1 = 2.38134142338928e-17 wuc1 = 9.24446373305873e-33 puc1 = 3.30607786168768e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.98 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.48333098191429+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.09657708623719e-07 wvth0 = 2.09602055374631e-07 pvth0 = -4.86786101463708e-14   k1 = -5.32540634376537 lk1 = 1.46493333415262e-06 wk1 = 2.29453179762791e-06 pk1 = -5.32888948276499e-13   k2 = 1.51733550138551 lk2 = -3.97808600727364e-07 wk2 = -5.51365528772814e-07 pk2 = 1.28050784498785e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 769244.314285716 lvsat = -0.150928295886657 wvsat = -0.233326970215677 pvsat = 5.41885555437995e-8   ua = -3.16602520721077e-09 lua = 1.69354477087854e-16 wua = 5.77048335283351e-16 pua = -1.34015436531211e-22   ub = 4.71931236044535e-18 lub = -6.09048897565707e-25 wub = -1.55661233942105e-24 pub = 3.61512319544163e-31   uc = 1.43601987732703e-13 luc = -1.58496608252677e-20 wuc = -3.06490088554054e-19 puc = 7.11801776360592e-26   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00432733337220327 lu0 = 1.5400672862666e-09 wu0 = 4.44485107156706e-09 pu0 = -1.03228554741395e-15   a0 = -12.2138655241736 la0 = 3.13866324103064e-06 wa0 = 8.79263718561222e-06 pa0 = -2.04202843789814e-12   keta = -0.44388971200618 lketa = 1.17112024060454e-07 wketa = 5.2946867553449e-07 pketa = -1.22965393612157e-13   a1 = 0.0   a2 = -8.88967409888088 la2 = 2.21984373557916e-06 wa2 = 4.25257907528117e-06 pa2 = -9.87631722180523e-13   ags = 24.2060879593981 lags = -5.3313907359545e-06 wags = -1.33226161506302e-05 pags = 3.09408434267081e-12   b0 = -7.14315972652866e-06 lb0 = 1.64255063062419e-12 wb0 = 3.60245672331625e-12 pb0 = -8.36645356793136e-19   b1 = -6.21689682938944e-07 lb1 = 1.44463442402509e-13 wb1 = 3.04586979482168e-13 pb1 = -7.07381938758772e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {7.82601577927585+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.86452850227436e-06 wvoff = -3.87316524915573e-06 pvoff = 8.99515516959674e-13   nfactor = {39.7759226071769+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -8.92514905096789e-06 wnfactor = -2.0603649696901e-05 pnfactor = 4.78505341655737e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -7.58075284287304 leta0 = 1.78929765420855e-06 weta0 = 3.59284951835771e-06 peta0 = -8.34414150691949e-13   etab = -1.58484448287688 letab = 3.45102919457446e-07 wetab = 4.75486749672683e-07 petab = -1.10428469204233e-13   dsub = 0.0600262179869873 ldsub = 4.66982431130687e-08 wdsub = 1.02237543178078e-07 pdsub = -2.37439537403065e-14   voffl = 0.0   minv = 0.0   pclm = 17.8463172396948 lpclm = -3.9993014554509e-06 wpclm = -8.41603091432391e-06 ppclm = 1.95456426763533e-12   pdiblc1 = 7.4195400363536 lpdiblc1 = -1.68385153661938e-06 wpdiblc1 = -3.58412693511157e-06 ppdiblc1 = 8.32388391791116e-13   pdiblc2 = 0.150326718036079 lpdiblc2 = -3.41269448100145e-08 wpdiblc2 = -7.28903137919829e-08 ppdiblc2 = 1.69282651459915e-14   pdiblcb = -2.48721704126105 lpdiblcb = 5.77637403882962e-07 wpdiblcb = 1.46751613954921e-06 ppdiblcb = -3.40820350797327e-13   drout = 1.0   pscbe1 = 801421942.103775 lpscbe1 = -0.330236100006914 wpscbe1 = -0.697252438862051 ppscbe1 = 1.61931998157727e-7   pscbe2 = -3.96943359392233e-08 lpscbe2 = 9.45097466153305e-15 wpscbe2 = -7.81915639458985e-15 ppscbe2 = 1.81594433854872e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 14.7195417797333 lbeta0 = -1.4731933109785e-06 wbeta0 = -1.07418442146732e-06 pbeta0 = 2.49471812594837e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.63973997086246e-08 lagidl = -2.7362587872542e-15 wagidl = 4.47687224593743e-15 pagidl = -1.03972224101324e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 2.44020055746748 lkt1 = -7.11313989867918e-07 wkt1 = -1.43649776382555e-06 pkt1 = 3.33616550164138e-13   kt2 = -0.12   at = 1073946.58415204 lat = -0.227310294345222 wat = -0.359177731420991 pat = 8.34165138784051e-8   ute = 6.86990560618665 lute = -1.62616911042761e-06 wute = -3.87016670129347e-06 pute = 8.988191252085e-13   ua1 = -7.58066301384651e-10 lua1 = 2.14498775822476e-16 wua1 = 5.00290881688466e-16 pua1 = -1.16189055235974e-22   ub1 = 5.34787479275022e-19 lub1 = -3.76576170292693e-26 wub1 = -7.95093731869616e-26 pub1 = 1.84654953570596e-32   uc1 = 7.46630777767922e-10 luc1 = -1.67751621961155e-16 wuc1 = -3.55191604668722e-16 puc1 = 8.2490763843078e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.99 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.026354617404+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -9.56080185470355e-10   k1 = 0.5362055478872 wk1 = -2.82146684111039e-8   k2 = -0.04000919904755 wk2 = 2.59757872776072e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -129809.6576462 wvsat = 0.075661676745305   ua = -1.3321200961346e-09 wua = 2.09577955309495e-16   ub = 1.1217330420374e-18 wub = -2.08960349801002e-25   uc = -1.957416097178e-11 wuc = -2.37504005485479e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.004827859608188 wu0 = 7.54683267220137e-10   a0 = 0.297555468698 wa0 = 4.67490181481865e-7   keta = -0.040513385789048 wketa = 2.34981636518712e-8   a1 = 0.0   a2 = 0.24699797 wa2 = 2.71165762014966e-7   ags = 0.5092246601128 wags = -1.34484788797876e-7   b0 = 1.3189463245e-08 wb0 = -4.93297414432489e-15   b1 = 8.49682495002e-09 wb1 = -3.0656451534772e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.3153511426394+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 5.30343278895116e-8   nfactor = {-0.921005428150001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.16308704081103e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0061742549595316 wpclm = -2.17423173621155e-9   pdiblc1 = 0.39   pdiblc2 = -0.0035349350792218 wpdiblc2 = 2.14421705723915e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 1191870692.5782 wpscbe1 = -197.010462048662   pscbe2 = 8.460328002298e-09 wpscbe2 = 5.18542742992053e-16   pvag = 0.0   delta = 0.01   alpha0 = 3.77194e-10 walpha0 = -1.359226877268e-16   alpha1 = 3.77194e-10 walpha1 = -1.359226877268e-16   beta0 = -71.84238 wbeta0 = 3.6699125686236e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.8619853383836e-09 wagidl = -8.28115689556303e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.0442122546 wkt1 = 2.5429775646807e-7   kt2 = -0.03455907535778 wkt2 = -8.78952623314677e-9   at = -197999.7942425 wat = 0.101993156706357   ute = -3.9171251944 wute = 1.30317236084947e-6   ua1 = -2.6829376059882e-09 wua1 = 1.19002967674905e-15   ub1 = 1.1853392376228e-18 wub1 = -3.38832996366663e-25   uc1 = -1.6084926039996e-10 wuc1 = 8.28912740197133e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.100 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08019591419462+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.07963876668072e-06 wvth0 = 2.54451181466652e-08 pvth0 = -5.29403244447179e-13   k1 = 0.555334390725375 lk1 = -3.83576204899898e-07 wk1 = -3.75945385802573e-08 pk1 = 1.88087435940317e-13   k2 = -0.063706997609727 lk2 = 4.75194015333824e-07 wk2 = 3.75960549377275e-08 pk2 = -2.33012430845774e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -201916.483938589 lvsat = 1.44590360277378 wvsat = 0.111019417652796 pvsat = -7.09002012608049e-7   ua = -1.36163064733859e-09 lua = 5.91752743806264e-16 wua = 2.24048519015582e-16 pua = -2.90167259781437e-22   ub = 1.23785605149496e-18 lub = -2.32852680353422e-24 wub = -2.65901522959135e-25 pub = 1.14179824087197e-30   uc = -1.1033584454605e-11 luc = -1.71257715682487e-16 wuc = -2.7938291033013e-17 puc = 8.39765976518821e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00538664936743245 lu0 = -1.12049880382809e-08 wu0 = 4.80679479437153e-10 pu0 = 5.49439053554476e-15   a0 = -0.311682338490566 la0 = 1.22165845545322e-05 wa0 = 7.66231280559953e-07 pa0 = -5.9904291128009e-12   keta = -0.0677749791532863 lketa = 5.46656094706894e-07 wketa = 3.68659459335309e-08 pketa = -2.68054018682934e-13   a1 = 0.0   a2 = -0.124077590421107 la2 = 7.44089730892523e-06 wa2 = 4.53123479433689e-07 pa2 = -3.64866036540557e-12   ags = 0.675130515746697 lags = -3.32678453229382e-06 wags = -2.1583709010084e-07 pags = 1.63129611433625e-12   b0 = 1.50492121126042e-08 lb0 = -3.72921362121748e-14 wb0 = -5.84490609300213e-15 pb0 = 1.82862810343396e-20   b1 = 8.66967920017286e-09 lb1 = -3.46611542764778e-15 wb1 = -3.150404615319e-15 pb1 = 1.69961732540103e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.379193158286858+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.28017561137262e-06 wvoff = 8.43394007146767e-08 pvoff = -6.27736927422907e-13   nfactor = {-1.78579990475459+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.73410689899331e-05 wnfactor = 1.58714091496194e-06 pnfactor = -8.50323132956547e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 6.99860641074996e-07 lcit = 1.86488654359028e-10 wcit = 4.56034379495546e-12 pcit = -9.14451219399892e-17   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 1.14599558634961 lpclm = -2.28559743136174e-05 wpclm = -5.61088129190266e-07 ppclm = 1.12074772878258e-11   pdiblc1 = 0.39   pdiblc2 = -0.00710017008226399 lpdiblc2 = 7.14909586331077e-08 wpdiblc2 = 3.89243788449789e-09 ppdiblc2 = -3.50557488458533e-14   pdiblcb = -0.225   drout = 0.56   pscbe1 = 1456711765.51736 lpscbe1 = -5310.65755095673 wpscbe1 = -326.875864814739 ppscbe1 = 0.00260409261355824   pscbe2 = 7.69142242655081e-09 lpscbe2 = 1.54182814489374e-14 wpscbe2 = 8.95577283651949e-16 ppscbe2 = -7.56038822870564e-21   pvag = 0.0   delta = 0.01   alpha0 = 5.631967871785e-10 lalpha0 = -3.72977308718057e-15 walpha0 = -2.27129563625909e-16 palpha0 = 1.82890243879978e-21   alpha1 = 5.631967871785e-10 lalpha1 = -3.72977308718057e-15 walpha1 = -2.27129563625909e-16 palpha1 = 1.82890243879978e-21   beta0 = -118.667338057552 lbeta0 = 0.000938945437434847 wbeta0 = 5.96598468846645e-05 pbeta0 = -4.6041396092614e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 3.38369940386337e-09 lagidl = -1.04615372175183e-14 wagidl = -1.08393932933525e-15 pagidl = 5.12983778999195e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.13721364818925 lkt1 = 1.86488654359028e-06 wkt1 = 2.99901194417625e-07 pkt1 = -9.14451219399892e-13   kt2 = -0.0345590753577801 wkt2 = -8.78952623314677e-9   at = -197999.7942425 wat = 0.101993156706357   ute = -3.9171251944 wute = 1.30317236084947e-6   ua1 = -2.6829376059882e-09 wua1 = 1.19002967674905e-15   ub1 = 1.1853392376228e-18 wub1 = -3.38832996366663e-25   uc1 = -1.73497449928098e-10 luc1 = 2.53624569928278e-16 wuc1 = 8.90933415808527e-17 puc1 = -1.24365365838385e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.101 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.966254849981498+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.62157629958033e-07 wvth0 = -3.39030816034583e-08 pvth0 = -5.15171184466472e-14   k1 = 0.56990211201905 lk1 = -5.00879036712839e-07 wk1 = -3.6651376143783e-08 pk1 = 1.80492862813352e-13   k2 = -0.0325947886498552 lk2 = 2.24670948522159e-07 wk2 = 2.00840593580163e-08 pk2 = -9.20015870230139e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -142577.639001077 lvsat = 0.968092803997611 wvsat = 0.0662930425442279 pvsat = -3.48854371724708e-7   ua = -1.53503300325172e-09 lua = 1.98803065039133e-15 wua = 2.82720809407433e-16 pua = -7.6261079938319e-22   ub = 1.23482799640303e-18 lub = -2.3041441681166e-24 wub = -2.28371973464514e-25 pub = 8.39601188660755e-31   uc = -1.4446517467789e-11 luc = -1.43775949717607e-16 wuc = -2.3943550950771e-17 puc = 5.18099797878291e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00314515910535934 lu0 = 6.84403623406533e-09 wu0 = 1.34055588252186e-09 pu0 = -1.42954321205923e-15   a0 = 1.21683434144772 la0 = -9.14031818840814e-08 wa0 = 1.81954288749211e-08 pa0 = 3.29373376789313e-14   keta = -0.0122351971917575 lketa = 9.94362741856475e-08 wketa = 8.02653578156043e-09 pketa = -3.58320801626013e-14   a1 = 0.0   a2 = 0.8   ags = 0.265503815399476 lags = -2.837080180981e-08 wags = -1.4517702013779e-08 pags = 1.0223480847929e-14   b0 = 8.85733456796954e-09 lb0 = 1.2566366403467e-14 wb0 = 5.02335742891139e-15 pb0 = -6.9227617832144e-20   b1 = 1.97010967519442e-08 lb1 = -9.22937701889759e-14 wb1 = -7.69316219487112e-15 pb1 = 3.82790052460465e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.259671906333613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.17761446980869e-07 wvoff = 2.28597199128715e-08 pvoff = -1.32687598044337e-13   nfactor = {-1.39843958725509+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.422194958487e-05 wnfactor = 1.17259526114182e-06 pnfactor = -5.16520899041196e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.38597e-05 wcit = -6.79613438634e-12   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -3.21364611818914 lpclm = 1.22489200842628e-05 wpclm = 1.37891822528936e-06 ppclm = -4.41392529998828e-12   pdiblc1 = 0.39   pdiblc2 = 0.0033367943719561 lpdiblc2 = -1.25500153346349e-08 wpdiblc2 = -1.02273599708054e-09 ppdiblc2 = 4.52242563586941e-15   pdiblcb = -0.225   drout = 0.56   pscbe1 = 759346316.573842 lpscbe1 = 304.698503740557 wpscbe1 = 10.1595909853236 ppscbe1 = -0.000109798776159619   pscbe2 = 9.3711305199161e-09 lpscbe2 = 1.89286371209358e-15 wpscbe2 = 4.13692541932535e-17 ppscbe2 = -6.82097602953085e-22   pvag = 0.0   delta = 0.01   alpha0 = 4.00796564076471e-10 lalpha0 = -2.42208702750882e-15 walpha0 = -1.08392703617397e-16 palpha0 = 8.72804388954263e-22   alpha1 = 4.82120308053189e-10 lalpha1 = -3.07692557567914e-15 walpha1 = -1.37697893671644e-16 palpha1 = 1.10877690043224e-21   beta0 = -81.0290838740599 lbeta0 = 0.0006358730686536 wbeta0 = 3.09379489344829e-05 pbeta0 = -2.29138259210076e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.1852827554532e-09 lagidl = -3.3020567149274e-14 wagidl = -1.92459903464924e-15 pagidl = 1.18990340174886e-20   bgidl = -229021220.317422 lbgidl = 9896.37751815242 wbgidl = 442.880500588068 pbgidl = -0.00356618141069677   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.46103623571751 lkt1 = 4.47238470725663e-06 wkt1 = 3.92788586377762e-07 pkt1 = -1.66240307109916e-12   kt2 = -0.00118574343781486 lkt2 = -2.68730178339216e-07 wkt2 = -2.21519821841788e-08 pkt2 = 1.07597742394505e-13   at = -459438.062529319 lat = 2.10516446574466 wat = 0.20396073674679 pat = -8.21067732607513e-7   ute = -8.32339191843367 lute = 3.54803303847331e-05 wute = 3.01887492308825e-06 pute = -1.38152539468693e-11   ua1 = -6.91302083941454e-09 lua1 = 3.40616581057746e-14 wua1 = 2.95092612392889e-15 pua1 = -1.41791660905288e-20   ub1 = 2.79014182596762e-18 lub1 = -1.29222604083815e-23 wub1 = -1.09047442770808e-24 pub1 = 6.0523994540289e-30   uc1 = 6.86213111740351e-12 luc1 = -1.19867460402829e-15 wuc1 = 2.67801250738914e-17 puc1 = 3.77395795587279e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.102 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.838274060758115+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.56451627306904e-07 wvth0 = -7.07775368618184e-08 pvth0 = 9.7907134752858e-14   k1 = 0.433111016898182 lk1 = 5.34317209530299e-08 wk1 = 2.08743095334689e-08 pk1 = -5.2615194292492e-14   k2 = 0.0628785977327022 lk2 = -1.62210413132855e-07 wk2 = -1.89470292954237e-08 pk2 = 6.61618687552679e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 210634.67662984 lvsat = -0.463209329531562 wvsat = -0.0639423634652967 pvsat = 1.78891140629546e-7   ua = -1.76376970045452e-09 lua = 2.91492733047449e-15 wua = 3.35580269941914e-16 pua = -9.76810178317817e-22   ub = 5.06676849516339e-19 lub = 6.46501219796946e-25 wub = 4.85232984721276e-26 pub = -2.82445738777599e-31   uc = -5.99617789449852e-11 luc = 4.06629499965312e-17 wuc = -9.38871110368901e-18 puc = -7.16976809862984e-24   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.000961403106718578 lu0 = 2.34848242120226e-08 wu0 = 3.04131005787463e-09 pu0 = -8.32141241385328e-15   a0 = 1.50606626539004 la0 = -1.26344122105587e-06 wa0 = -8.32094366930922e-08 pa0 = 4.43854494342854e-13   keta = 0.0519252828146405 lketa = -1.60557581796919e-07 wketa = -1.22221351371234e-08 pketa = 4.62204548269387e-14   a1 = 0.0   a2 = 0.8   ags = -0.639516382743009 lags = 3.63899096097169e-06 wags = 2.589364675808e-07 pags = -1.09787926371252e-12   b0 = 1.25088617165385e-07 lb0 = -4.58431034882934e-13 wb0 = -5.18897795826239e-14 pb0 = 1.61398243230891e-19   b1 = 1.57663276030461e-08 lb1 = -7.63491294487374e-14 wb1 = -7.53172723557841e-15 pb1 = 3.76248315622974e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0716933548956766+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.43973322233649e-07 wvoff = -4.95996044420371e-08 pvoff = 1.60935191857571e-13   nfactor = {1.94471644241471+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.7466896573271e-07 wnfactor = -4.09112082986595e-08 pnfactor = -2.47785894167059e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.38597e-05 wcit = -6.79613438634e-12   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.16157665925 leta0 = -3.30568446409198e-7   etab = -0.14131544425 letab = 2.88987509753953e-7   dsub = 0.86783645 ldsub = -1.24742809965735e-6   voffl = 0.0   minv = 0.0   pclm = 0.145058441069095 lpclm = -1.36136695505946e-06 wpclm = 1.74821619234141e-07 ppclm = 4.65366743222723e-13   pdiblc1 = 0.39   pdiblc2 = 0.00299154118364688 lpdiblc2 = -1.11509655190811e-08 wpdiblc2 = -1.18506076822936e-09 ppdiblc2 = 5.18020505348384e-15   pdiblcb = -0.999093746142 lpdiblcb = 3.1368159641477e-06 wpdiblcb = 2.78946384428511e-07 ppdiblcb = -1.13035853367574e-12   drout = 0.56   pscbe1 = 869979949.826348 lpscbe1 = -143.615862171473 wpscbe1 = -34.3148223532394 ppscbe1 = 7.04223539706788e-5   pscbe2 = 9.93818823893751e-09 lpscbe2 = -4.04991960406971e-16 wpscbe2 = -1.50234201441378e-16 ppscbe2 = 9.43261589181696e-23   pvag = 0.0   delta = 0.01   alpha0 = -4.13359598025765e-10 lalpha0 = 8.77071581276836e-16 walpha0 = 2.2196677453893e-16 palpha0 = -4.65892493888369e-22   alpha1 = -5.61626499026106e-10 lalpha1 = 1.15259011708029e-15 walpha1 = 2.75395078501585e-16 palpha1 = -5.65176204405921e-22   beta0 = 227.480776093434 lbeta0 = -0.000614283851830657 wbeta0 = -8.95428480008289e-05 pbeta0 = 2.59079206805463e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -3.32411957975479e-09 lagidl = 5.51384189775621e-15 wagidl = 1.55224995622615e-15 pagidl = -2.19000296784327e-21   bgidl = 3458042440.63485 lbgidl = -5044.50039249578 wbgidl = -885.761001176136 pbgidl = 0.00181779681433672   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.121060842409585 lkt1 = -9.57521200447667e-07 wkt1 = -8.41149537648774e-08 pkt1 = 2.70125961119067e-13   kt2 = -0.0714778799357591 lkt2 = 1.61106397396231e-08 wkt2 = 5.83332049092885e-09 pkt2 = -5.80550447358059e-15   at = 178112.277467314 lat = -0.478344436654314 wat = -0.0450370316086666 pat = 1.87931731226507e-7   ute = 2.29773887766882 lute = -7.55907253585768e-06 wute = -1.00242748573269e-06 pute = 2.48004059015852e-12   ua1 = 2.97725345581748e-09 lua1 = -6.01613667515929e-15 wua1 = -1.08315923988644e-15 pua1 = 2.16792808639434e-21   ub1 = -7.58384781229336e-19 lub1 = 1.45723169594614e-24 wub1 = 5.32704661397096e-25 pub1 = -5.25116647543923e-31   uc1 = -6.39347534736526e-10 luc1 = 1.41992399096063e-15 wuc1 = 2.46181708237271e-16 puc1 = -5.11672733975443e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.103 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.13425382143309+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.5097076467999e-07 wvth0 = 1.1125377856542e-08 pvth0 = -7.0177548657495e-14   k1 = 0.31600760780741 lk1 = 2.93756372535703e-07 wk1 = 4.70912272089895e-08 pk1 = -1.06418680073655e-13   k2 = -0.00729958632938632 lk2 = -1.81877261387223e-08 wk2 = 7.57891917199489e-09 pk2 = 1.17241766946473e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -229978.447576143 lvsat = 0.441035870328296 wvsat = 0.100780667432531 pvsat = -1.59160546469304e-7   ua = 2.31929699434257e-09 lua = -5.46451771245597e-15 wua = -9.21408826400807e-16 pua = 1.60283689572786e-21   ub = -7.68265742368126e-19 lub = 3.26299322939369e-24 wub = 3.79014321976481e-25 pub = -9.60693628327244e-31   uc = -1.12789601842919e-10 luc = 1.49078479744055e-16 wuc = 1.38964357577427e-18 puc = -2.92895710410757e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.021315975733608 lu0 = -2.22337705713858e-08 wu0 = -4.11453164128967e-09 pu0 = 6.36411362236477e-15   a0 = -0.314983504150515 la0 = 2.47379542113535e-06 wa0 = 6.93392247852833e-07 pa0 = -1.14992087655473e-12   keta = -0.0794469659022819 lketa = 1.09050196026644e-07 wketa = 3.3312058277737e-08 pketa = -4.72267748693544e-14   a1 = 0.0   a2 = 2.387598984568 la2 = -3.25813890288679e-06 wa2 = -5.72094786806845e-07 pa2 = 1.17407752156084e-12   ags = 2.38711338853533 lags = -2.57238880072589e-06 wags = -8.29264887373017e-07 pags = 1.13537434958197e-12   b0 = -2.47448155666944e-07 lb0 = 3.06104949404805e-13 wb0 = 5.06499908600982e-14 pb0 = -4.90382828817924e-20   b1 = -2.9174994021583e-08 lb1 = 1.58813832661562e-14 wb1 = 9.40017166061047e-15 pb1 = 2.87646057588601e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.431578643362545+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.94598741825463e-07 wvoff = 7.80493084165309e-08 pvoff = -1.01031396014035e-13   nfactor = {3.09192789495963+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.67968770727242e-06 wnfactor = -2.73812456433529e-07 pnfactor = 2.3018406200899e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.38597e-05 wcit = -6.79613438634e-12   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.5145729485 leta0 = 1.05705485304849e-06 weta0 = 2.81241408268029e-23 peta0 = -9.19022954582479e-29   etab = -0.0680382695671501 letab = 1.38604940951297e-07 wetab = 1.17994549778912e-07 petab = -2.42153488821923e-13   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = -1.91213007960055 lpclm = 2.86048378616518e-06 wpclm = 8.90306993711852e-07 ppclm = -1.00298310815154e-12   pdiblc1 = 0.378118783024182 lpdiblc1 = 2.43831443701047e-08 wpdiblc1 = 5.56363610406627e-09 ppdiblc1 = -1.14179332491172e-14   pdiblc2 = -0.00546406055573012 lpdiblc2 = 6.20198396134312e-09 wpdiblc2 = 2.74817238731051e-09 ppdiblc2 = -2.89174515734077e-15   pdiblcb = 1.323187492284 lpdiblcb = -1.62906945144339e-06 wpdiblcb = -5.57892768857023e-07 ppdiblcb = 5.8703876078042e-13   drout = -0.213856349057381 ldrout = 1.58814127535857e-06 wdrout = 2.10033130475658e-07 pdrout = -4.31039021786756e-13   pscbe1 = 735932637.192775 lpscbe1 = 131.48179684959 wpscbe1 = 32.0366501521785 ppscbe1 = -6.57469910182572e-5   pscbe2 = 1.06266885376439e-08 lpscbe2 = -1.81796187892507e-15 wpscbe2 = -2.70009306685044e-16 ppscbe2 = 3.40133780228744e-22   pvag = 0.0   delta = 0.01   alpha0 = -7.64670602543543e-11 lalpha0 = 1.85686228883223e-16 walpha0 = -1.03627346082709e-17 palpha0 = 1.09041149524108e-23   alpha1 = -1.05228234160545e-10 lalpha1 = 2.15949972797794e-16 walpha1 = 1.41768340749623e-21 palpha1 = -1.49174744175405e-27   beta0 = -160.356629202232 lbeta0 = 0.000181652748325536 wbeta0 = 7.75613634048155e-05 pbeta0 = -8.38592413222906e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.57207713019799e-10 lagidl = -2.24636056954939e-15 wagidl = -1.95066518947785e-16 pagidl = 1.39591503711712e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.577486688374741 lkt1 = -2.0824453046599e-08 wkt1 = 5.6928802500759e-08 pkt1 = -1.93301003707917e-14   kt2 = -0.0767464696527841 lkt2 = 2.69230661062595e-08 wkt2 = 1.05825485297624e-08 pkt2 = -1.55520744716806e-14   at = -227146.005284984 lat = 0.35334403731611 wat = 0.114003357437388 pat = -1.38457793910536e-7   ute = -4.25228135467153 lute = 5.88316063582119e-06 wute = 1.20664662991352e-06 pute = -2.05351630015761e-12   ua1 = -4.25727796880758e-09 lua1 = 8.83087979930752e-15 wua1 = 1.56101111156054e-15 pua1 = -3.25855200817025e-21   ub1 = 4.23303914067593e-18 lub1 = -8.78638310781648e-24 wub1 = -1.30512493951958e-24 pub1 = 3.24655628613011e-30   uc1 = 1.98840461012325e-10 luc1 = -3.00241455998979e-16 wuc1 = -4.97368913523963e-17 puc1 = 9.56241406022539e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.104 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.869619937697598+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.74883870434939e-08 wvth0 = -6.56968270884723e-08 pvth0 = 1.06580787404616e-14   k1 = 0.583519059636835 lk1 = 1.22693199283541e-08 wk1 = -7.63322974537229e-08 pk1 = 2.34528597880112e-14   k2 = -0.00196952681590132 lk2 = -2.37962439513703e-08 wk2 = 2.19166294983317e-08 pk2 = -3.36257863226827e-15   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 346531.375966435 lvsat = -0.165592555925616 wvsat = -0.118709456039089 pvsat = 7.17963995228433e-8   ua = -3.44757910171813e-09 lua = 6.0363729149123e-16 wua = 9.5887270804047e-16 pua = -3.75676186917235e-22   ub = 2.6019529638409e-18 lub = -2.83295812683812e-25 wub = -7.92049779575943e-25 pub = 2.71550375082584e-31   uc = 4.74258562501869e-11 luc = -1.95071145262091e-17 wuc = -4.20119614100521e-17 puc = 1.63794639940253e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00282560961218074 lu0 = 3.16904361762304e-09 wu0 = 3.34242424654504e-09 pu0 = -1.48241601191809e-15   a0 = 3.43911487494707 la0 = -1.47642831958143e-06 wa0 = -1.02398735509863e-06 pa0 = 6.57179788993727e-13   keta = -0.0119187782793133 lketa = 3.79941332976888e-08 wketa = 1.14382589939114e-08 pketa = -2.42102226895439e-14   a1 = 0.0   a2 = -2.375197969136 la2 = 1.75348085206957e-06 wa2 = 1.14418957361369e-06 pa2 = -6.31870682701145e-13   ags = 0.202869707650952 lags = -2.74033677221067e-07 wags = -8.47185484005195e-08 pags = 3.51930676222531e-13   b0 = 3.64226845093589e-07 lb0 = -3.3752578842046e-13 wb0 = -8.72699363082923e-14 pb0 = 9.60869950416564e-20   b1 = -2.25641708810144e-08 lb1 = 8.9251908922549e-15 wb1 = 2.2161307974218e-14 pb1 = -1.05513557821533e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.105472179516606+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.85445020111791e-08 wvoff = -3.35774299771274e-08 pvoff = 1.64270580735231e-14   nfactor = {1.19460064249209+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.16761612845773e-07 wnfactor = -1.71154584027989e-07 pnfactor = 1.22163034375367e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 3.91675446142e-05 lcit = -1.61075723403797e-11 wcit = -1.43023696701711e-11 pcit = 7.89838353376431e-18   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 0.134040766574684 letab = -7.4031310275695e-08 wetab = -2.35993790954876e-07 petab = 1.3032826479682e-13   dsub = 0.338527019695156 ldsub = -8.26295067850904e-08 wdsub = -5.88954232839957e-08 pdsub = 6.19722968826215e-14   voffl = 0.0   minv = 0.0   pclm = 1.0777156784583 lpclm = -2.85560483831945e-07 wpclm = -1.70285638329201e-07 ppclm = 1.13018064765236e-13   pdiblc1 = 1.10211910979743 lpdiblc1 = -7.37441131474759e-07 wpdiblc1 = -2.43690347837194e-07 ppdiblc1 = 2.50857826575186e-13   pdiblc2 = 0.00260978353966874 lpdiblc2 = -2.29366197113165e-09 wpdiblc2 = -1.34316012702475e-09 ppdiblc2 = 1.4133308415409e-15   pdiblcb = 0.387313784568 lpdiblcb = -6.44302893615186e-07 wpdiblcb = -3.00249411353245e-07 ppdiblcb = 3.15935341350573e-13   drout = 1.87425700408743 ldrout = -6.09061383694589e-07 wdrout = -4.54736615941685e-07 pdrout = 2.6846029049267e-13   pscbe1 = 928134725.61445 lpscbe1 = -70.7615052775013 wpscbe1 = -64.073300304357 ppscbe1 = 3.53840315799791e-5   pscbe2 = 4.30053949738211e-08 lpscbe2 = -3.58882290754474e-14 wpscbe2 = -1.23341256806818e-14 ppscbe2 = 1.30345157859522e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 16.578854573318 lbeta0 = -4.52637592889996e-06 wbeta0 = -4.85803889610213e-06 pbeta0 = 2.86599781303381e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.86785712268797e-09 lagidl = 1.25241562837026e-15 wagidl = 1.87848672609837e-15 pagidl = -7.85966850109987e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.694336388564203 lkt1 = 1.02129826029861e-07 wkt1 = 8.11456671180289e-08 pkt1 = -4.48121266462617e-14   kt2 = -0.0912884341855341 lkt2 = 4.2224746492094e-08 wkt2 = 2.40800167543872e-08 pkt2 = -2.97546909287644e-14   at = 115957.061969135 lat = -0.00768376348056543 wat = -0.0174223577679177 pat = -1.66005065759252e-10   ute = 2.76184731451803 lute = -1.49740715743285e-06 wute = -1.49055761187952e-06 pute = 7.84597982839427e-13   ua1 = 8.60599439777334e-09 lua1 = -4.70440850552069e-15 wua1 = -3.35392428463804e-15 pua1 = 1.91315435793193e-21   ub1 = -9.23566631966808e-18 lub1 = 5.38596793189228e-24 wub1 = 3.76829351605467e-24 pub1 = -2.0919127698187e-30   uc1 = -2.08887045083974e-10 luc1 = 1.28786958198309e-16 wuc1 = 8.65776896698688e-17 puc1 = -4.78119230763574e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.105 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.839540480836513+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.40995565388301e-08 wvth0 = -1.0249013656543e-07 pvth0 = 3.09769263459452e-14   k1 = 0.636553775766274 lk1 = -1.70187308111162e-08 wk1 = -7.48044686188999e-08 pk1 = 2.26091270087822e-14   k2 = -0.0691573633633802 lk2 = 1.33077684671191e-08 wk2 = 3.49629063671156e-08 pk2 = -1.05672937091161e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -4003.15547101782 lvsat = 0.0279876853189968 wvsat = 0.0249597335657953 pvsat = -7.54390475212666e-9   ua = -3.39394382705758e-09 lua = 5.74017586506866e-16 wua = 6.15418215956633e-16 pua = -1.86005847845381e-22   ub = 2.92414273629912e-18 lub = -4.61222859195454e-25 wub = -6.63414285359095e-25 pub = 2.00512323849789e-31   uc = 2.66669143135392e-11 luc = -8.04313415428898e-18 wuc = -2.72853904437847e-17 puc = 8.24681826390081e-24   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.000880803098414026 lu0 = 1.12220314308605e-09 wu0 = 1.45365752506674e-09 pu0 = -4.39357811348745e-16   a0 = 0.70937693429585 la0 = 3.1050349977619e-08 wa0 = 3.66759760207981e-07 pa0 = -1.10850570204541e-13   keta = 0.137701308077867 lketa = -4.46325120524596e-08 wketa = -7.15740969118774e-08 pketa = 2.16327697729366e-14   a1 = 0.0   a2 = 1.13401084291128 la2 = -1.84455149921854e-7   ags = -1.15794989857545 lags = 4.77469424580219e-07 wags = 1.22058180359273e-06 pags = -3.68912306063278e-13   b0 = -5.45536251221767e-07 lb0 = 1.64884513178021e-13 wb0 = 1.91571134419824e-13 pb0 = -5.7901034380451e-20   b1 = -1.41428581103565e-08 lb1 = 4.2745798638485e-15 wb1 = 6.74828566981099e-15 pb1 = -2.03962210570069e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.186094070486154+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.02162707648335e-09 wvoff = -8.46337035734288e-09 pvoff = 2.55799444691443e-15   nfactor = {1.18995440327013+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.19327465932427e-07 wnfactor = 1.10576453711995e-07 pnfactor = -3.34209590992747e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 4.261986923225e-05 letab = -3.17717446363629e-11 wetab = 9.38279410478891e-12 petab = -2.83588383861372e-18   dsub = -0.341956085992193 ldsub = 2.93162524949008e-07 wdsub = 1.17790846567992e-07 pdsub = -3.56014588392495e-14   voffl = 0.0   minv = 0.0   pclm = 0.468101347119457 lpclm = 5.10947633496139e-08 wpclm = 7.59160519896122e-08 ppclm = -2.29450953014963e-14   pdiblc1 = -1.07369926187291 lpdiblc1 = 4.64139333551583e-07 wpdiblc1 = 4.65126151258122e-07 ppdiblc1 = -1.40581123334709e-13   pdiblc2 = -0.0167899269371855 lpdiblc2 = 8.41969234173775e-09 wpdiblc2 = 2.6863202540495e-09 ppdiblc2 = -8.11921492544683e-16   pdiblcb = -1.449627569136 lpdiblcb = 3.70135110378372e-07 wpdiblcb = 6.0049882270649e-07 ppdiblcb = -1.81496565671278e-13   drout = 1.18204717077318 ldrout = -2.26793348715629e-07 wdrout = 6.93407099807406e-08 pdrout = -2.0957744206709e-14   pscbe1 = 800086006.26808 lpscbe1 = -0.0474963595033842   pscbe2 = -5.96894384119651e-08 lpscbe2 = 2.08242737980193e-14 wpscbe2 = 2.48923248707018e-14 ppscbe2 = -7.52353094589551e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.28154809139276 lbeta0 = 6.07996494597877e-07 wbeta0 = 7.32719355734711e-07 pbeta0 = -2.21459296235328e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.44625077053725e-09 lagidl = 4.67343471639489e-16 wagidl = 1.00565717988303e-15 pagidl = -3.03952843019386e-22   bgidl = 664683394.7904 lbgidl = 185.176248010765   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.50617204476 lkt1 = -1.78261568560336e-9   kt2 = -0.0114863736473116 lkt2 = -1.84538282571557e-09 wkt2 = -6.58266809450854e-08 pkt2 = 1.98956535288855e-14   at = 144946.508737821 lat = -0.0236929825324454 wat = -0.0391495207463496 pat = 1.1832668598939e-8   ute = 0.335200998754125 lute = -1.57308716076443e-07 wute = -1.54208097671027e-07 pute = 4.66083180643841e-14   ua1 = -2.93892954124587e-10 lua1 = 2.10491985353478e-16 wua1 = 2.43892596842241e-16 pua1 = -7.37148301473895e-23   ub1 = 6.11804718079272e-19 lub1 = -5.22290164064338e-26 wub1 = -4.3596214528491e-26 pub1 = 1.31766506677348e-32   uc1 = 5.303025600552e-11 luc1 = -1.58550379072564e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.106 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.900132306847143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.57861012698991e-8   k1 = -0.753854237424425 lk1 = 4.03222358319681e-7   k2 = 0.540335591016728 lk2 = -1.70907210543588e-07 pk2 = -1.89326617253043e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -13507.8828004287 lvsat = 0.0308604226212199   ua = 1.63077910708429e-09 lua = -9.44669747276976e-16   ub = -9.19993558705713e-19 lub = 7.00640427015691e-25   uc = -1.06695290525572e-14 luc = 1.99788190474911e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0121906473150571 lu0 = -2.29611810248482e-9   a0 = -0.80891296242857 la0 = 4.89942843233298e-7   keta = -0.243357161001197 lketa = 7.0539742817404e-08 wketa = -1.98523347012727e-23 pketa = 4.73316543132607e-30   a1 = 0.0   a2 = 0.0430362205630015 la2 = 1.45284292860557e-7   ags = -2.32595109449885 lags = 8.30489610039697e-07 pags = 1.0097419586829e-28   b0 = 2.34260196342857e-07 lb0 = -7.08035045232542e-14   b1 = -1.14807668171428e-09 lb1 = 3.46998140511371e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.189659108206143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.94411938088082e-9   nfactor = {5.23503302213285+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.03269231068501e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.70540283255443 leta0 = -3.67346998319748e-7   etab = 0.327817537026143 letab = -9.90994460308925e-08 wetab = 1.96455395481344e-23 petab = 9.83610941197449e-30   dsub = 1.84528256562071 ldsub = -3.67915046830431e-07 pdsub = 1.0097419586829e-28   voffl = 0.0   minv = 0.0   pclm = 0.674204565135856 lpclm = -1.11984915733169e-8   pdiblc1 = 1.43337925002629 lpdiblc1 = -2.93607597120365e-7   pdiblc2 = 0.0365667326803343 lpdiblc2 = -7.70698453104027e-9   pdiblcb = -0.971476165276739 lpdiblcb = 2.25617195621737e-7   drout = -1.453869509709 ldrout = 5.69894016543347e-7   pscbe1 = 799692834.756857 lpscbe1 = 0.0713369775635329   pscbe2 = 3.64473694867385e-08 lpscbe2 = -8.23240343170863e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 12.33537434018 lbeta0 = -9.19487112314327e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.48814030467986e-08 lagidl = 4.52802420107354e-15 wagidl = 1.08468374467889e-30 pagidl = -2.82118644197349e-37   bgidl = 2197559304.32 lbgidl = -278.124765513191   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.145358303 lkt1 = -1.10836043436371e-7   kt2 = 0.322172873485714 lkt2 = -1.02691554656943e-07 wkt2 = -2.64697796016969e-23 pkt2 = 6.31088724176809e-30   at = -28431.3870000001 lat = 0.028709272809041   ute = -0.361641969714286 lute = 5.33071932423549e-8   ua1 = 1.18888162042857e-09 lua1 = -2.37666250383193e-16   ub1 = 6.59166363999999e-19 lub1 = -6.65437423544519e-26   uc1 = -7.82166285911428e-11 luc1 = 2.38134142338928e-17 wuc1 = 3.08148791101958e-33 puc1 = 1.0101904577379e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.107 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -2.61215e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.98239e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.384395e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.52479736550476+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.19287985947923e-07 wvth0 = 2.2993518779427e-07 pvth0 = -5.34008378189046e-14   k1 = -4.31069232248112 lk1 = 1.2292731057075e-06 wk1 = 1.79696454492033e-06 pk1 = -4.17332436805932e-13   k2 = 1.39494703504205 lk2 = -3.69384736138362e-07 wk2 = -4.91352075046678e-07 pk2 = 1.14113079965066e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 886155.684141414 lvsat = -0.178080143156054 wvsat = -0.290654717629433 pvsat = 6.75025235864124e-8   ua = -1.05119578754181e-09 lua = -3.21799851824331e-16 wua = -4.59962923276053e-16 pua = 1.068231691904e-22   ub = 1.71549560447035e-18 lub = 8.85665172921955e-26 wub = -8.36841847318501e-26 pub = 1.94350661146787e-32   uc = 7.84407846329833e-13 luc = -1.64672335843441e-19 wuc = -6.20710651090046e-19 puc = 1.44155703741106e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0121002679748236 lu0 = -2.27512813337096e-09 wu0 = -3.61045938967053e-09 pu0 = 8.38503920035252e-16   a0 = 9.92751868810672 la0 = -2.00351825258197e-06 wa0 = -2.06443927392469e-06 pa0 = 4.79451570294092e-13   keta = 1.33334916229022 lketa = -2.95639263822766e-07 wketa = -3.42004316402275e-07 pketa = 7.94281084542135e-14   a1 = 0.0   a2 = -5.03122926223924 la2 = 1.323746931383e-06 wa2 = 2.36058216105529e-06 pa2 = -5.48228682829964e-13   ags = -14.6426762795833 lags = 3.69096281719928e-06 wags = 5.72696086123568e-06 pags = -1.33004657129596e-12   b0 = 1.06228498170058e-06 lb0 = -2.63106464749089e-13 wb0 = -4.21101141342315e-13 pb0 = 9.77977923687632e-20   b1 = -3.1811861423236e-08 lb1 = 7.46844750023661e-15 wb1 = 1.53390919707336e-14 pb1 = -3.56239673655909e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.418287926502107+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 5.0153323266629e-08 wvoff = 1.69447210440644e-07 pvoff = -3.93529284943665e-14   nfactor = {-6.80141393539786+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.89211131968931e-06 wnfactor = 2.23564974689098e-06 pnfactor = -5.19214004167201e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -2.17198988115483 leta0 = 5.33150317690232e-07 weta0 = 9.4065070080067e-07 peta0 = -2.1845954070605e-13   etab = -1.06884986240379 letab = 2.25266780814914e-07 wetab = 2.22467652335536e-07 petab = -5.16665549813619e-14   dsub = 0.268524401900667 ldsub = -1.72400061359654e-9   voffl = 0.0   minv = 0.0   pclm = 3.85946465030683 lpclm = -7.50952849533679e-07 wpclm = -1.55754697604184e-06 ppclm = 3.61729382356884e-13   pdiblc1 = 2.72941641280929 lpdiblc1 = -5.94603155916578e-07 wpdiblc1 = -1.28431449803465e-06 ppdiblc1 = 2.9827305196706e-13   pdiblc2 = 0.0624245614186734 lpdiblc2 = -1.37122842507184e-08 wpdiblc2 = -2.97872979098934e-08 ppdiblc2 = 6.91789142848738e-15   pdiblcb = 1.90433904108104 lpdiblcb = -4.42270755348411e-07 wpdiblcb = -6.85893046850613e-07 ppdiblcb = 1.59293858879727e-13   drout = -0.687671721436047 ldrout = 3.91949943601472e-07 wdrout = 8.27553541483953e-07 pdrout = -1.92193517134858e-13   pscbe1 = 744593680.431477 lpscbe1 = 12.8677298755529 wpscbe1 = 27.1686106943271 ppscbe1 = -6.30971965348299e-6   pscbe2 = -8.00542949772542e-08 lpscbe2 = 1.88242926284024e-14 wpscbe2 = 1.19714383116185e-14 ppscbe2 = -2.78028274780521e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 30.6038043877617 lbeta0 = -5.16220211185483e-06 wbeta0 = -8.86306753669177e-06 pbeta0 = 2.05838539392391e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 3.22217720971693e-08 lagidl = -6.41135850388697e-15 wagidl = -3.28264356840471e-15 pagidl = 7.62370990257015e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.119882863924222 lkt1 = -1.16752535833647e-07 wkt1 = -1.81155225962607e-07 pkt1 = 4.20720331432335e-14   kt2 = -0.12   at = 447224.86482124 lat = -0.0817585620826792 wat = -0.0518633575593503 pat = 1.20449017496562e-8   ute = -4.05204580269321 lute = 9.10377650624879e-07 wute = 1.48543620034386e-06 pute = -3.4498215947646e-13   ua1 = -1.274186416869e-10 lua1 = 6.80352713912908e-17 wua1 = 1.91051414330822e-16 pua1 = -4.43703536184331e-23   ub1 = 3.7264e-19   uc1 = 2.72225892665131e-10 luc1 = -5.7574408230228e-17 wuc1 = -1.22566125567821e-16 puc1 = 2.84651247002475e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.07365e-11   cgso = 6.07365e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.10485215e-11   cgdl = 1.10485215e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -1.51275e-8   dwc = 2.252e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000787089375   mjs = 0.34629   pbs = 0.6587   cjsws = 1.05469e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.5506845e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__pfet_01v8





















