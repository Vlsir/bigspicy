** Translated using xdm 2.6.0 on Nov_14_2022_16_05_27_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__esd_pfet_g5v0d10v5 d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__esd_pfet_g5v0d10v5 d g s b sky130_fd_pr__esd_pfet_g5v0d10v5__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.0 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.4495e-05 wmax = 1.4505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.0072+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {154260+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.0216+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.55852+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0}   kt2 = 0.01   at = 0.0   ute = -1.115   ua1 = 1.56e-9   ub1 = -3.963e-18   uc1 = -8.9645e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.1 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.5495e-05 wmax = 1.5505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.0152+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {155260+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.021700+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.548+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1}   kt2 = 0.02   at = 0.0   ute = -1.121   ua1 = 5.4616e-10   ub1 = -2.0736e-18   uc1 = -2.000e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.2 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.6495e-05 wmax = 1.6505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.01918+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {152260+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.0219+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.548+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2}   kt2 = 0.02   at = 0.0   ute = -1.0681   ua1 = 8.227e-10   ub1 = -1.9492e-18   uc1 = -1.36e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.3 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.7495e-05 wmax = 1.7505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.01218+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {159860+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.02165+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.548+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3}   kt2 = 0.02   at = 0.0   ute = -1.0881   ua1 = 5.9616e-10   ub1 = -2.0036e-18   uc1 = -2.0e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.4 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.9495e-05 wmax = 1.9505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.01018+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {148260+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.022+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.538+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4}   kt2 = 0.02   at = 0.0   ute = -1.111   ua1 = 5.9616e-10   ub1 = -2.0736e-18   uc1 = -1.12e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.5 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 2.1495e-05 wmax = 2.1505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.01218+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {150260+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.0219+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.538+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5}   kt2 = 0.02   at = 0.0   ute = -1.115   ua1 = 5.9616e-10   ub1 = -2.0736e-18   uc1 = -1.3393e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.6 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 2.3495e-05 wmax = 2.3505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.01518+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {149560+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.022046+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.538+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6}   kt2 = 0.02   at = 0.0   ute = -1.095   ua1 = 8.3462e-10   ub1 = -2.0736e-18   uc1 = -1.0304e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* .model sky130_fd_pr__esd_pfet_g5v0d10v5__model.7 pmos  lmin = 5.45e-07 lmax = 5.55e-07 wmin = 2.6495e-05 wmax = 2.6505e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.175e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {1e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.53e-8   dwb = -1.0e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 200000.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.577   rnoib = 0.37   tnoia = 1.5   tnoib = 3.5   epsrox = 3.9   toxe = {1.175e-008*sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult}   vth0 = {-1.0172+sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7}   k1 = 0.64397   k2 = {0.0012758+sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7}   k3 = -1.584   dvt0 = 4.0   dvt1 = 0.39618   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-9   k3b = 0.24   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {150260+sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7}   ua = {2.718e-009+sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7}   ub = {1.5031e-018+sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7}   uc = 2.5114e-11   rdsw = {329.4+sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.022046+sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7}   a0 = {0.71809+sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7}   keta = {-0.01188+sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7}   a1 = 0.0   a2 = 0.5   ags = {0.097232+sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7}   b0 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7}   b1 = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15351+sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7}   nfactor = {1.1792+sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7}   cit = 1.0e-5   cdsc = 1.0e-5   cdscb = -0.00030725687   cdscd = 7.8783957e-11   eta0 = {0.0154+sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7}   etab = -6.956e-5   dsub = 0.10478   voffl = 0.0   minv = 0.0   pclm = {0.46878+sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7}   pdiblc1 = 0.0   pdiblc2 = 0.0   pdiblcb = -0.5   drout = 0.46464   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.561e-6   alpha1 = 1.0e-10   beta0 = 36.0   fprout = 10.125   pdits = {1.1249e-012+sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7}   agidl = {7.25e-010+sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7}   bgidl = {1.334e+009+sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7}   cgidl = {650+sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7}   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.175e-8   kt1 = {-0.538+sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7}   kt2 = -0.02   at = 0.0   ute = -1.271   ua1 = 1.0114e-9   ub1 = -4.3718e-18   uc1 = -5.152e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0000000e+40   noib = 8.5300000e+24   noic = 8.4000000e+7   em = 4.1000000e+7   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 4.02e-12   xtis = 10.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.00096   tcjsw = 3.0e-5   tcjswg = 0.0   cgdo = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgso = {1.9771e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cgdl = {1.0005e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult}   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = {4.4983e-008+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak}   dwc = {0+sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff}   vfbcv = -0.1446893   acde = 0.401   moin = 15.773   noff = 4.0   voffcv = 0.0   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.00077547*sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult}   mjs = 0.33956   pbs = 0.6587   cjsws = {9.8717e-011*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjsws = 0.24676   pbsws = 1.0   cjswgs = {1.46e-010*sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult}   mjswgs = 0.81   pbswgs = 3.0; HSpice Parser Retained (as a comment). Continuing.










* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























.ENDS sky130_fd_pr__esd_pfet_g5v0d10v5










