** Translated using xdm 2.6.0 on Nov_14_2022_16_05_17_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 3
.PARAM 
+ SKY130_FD_PR__ESD_NFET_01V8__TOXE_MULT=1.052 SKY130_FD_PR__ESD_NFET_01V8__RSHN_MULT=1.0 
+ SKY130_FD_PR__ESD_NFET_01V8__OVERLAP_MULT=1.0257 SKY130_FD_PR__ESD_NFET_01V8__AJUNCTION_MULT=1.2169e+0 
+ SKY130_FD_PR__ESD_NFET_01V8__PJUNCTION_MULT=1.2474e+0 SKY130_FD_PR__ESD_NFET_01V8__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__ESD_NFET_01V8__WINT_DIFF=3.2175e-8 SKY130_FD_PR__ESD_NFET_01V8__DLC_DIFF=-14.422e-9 
+ SKY130_FD_PR__ESD_NFET_01V8__DWC_DIFF=3.2175e-8 SKY130_FD_PR__ESD_NFET_01V8__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__UA_DIFF_0=1.3831e-10 SKY130_FD_PR__ESD_NFET_01V8__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITSD_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__K2_DIFF_0=0.0017582 SKY130_FD_PR__ESD_NFET_01V8__UB_DIFF_0=-7.8945e-20 
+ SKY130_FD_PR__ESD_NFET_01V8__VTH0_DIFF_0=0.062077 SKY130_FD_PR__ESD_NFET_01V8__U0_DIFF_0=0.0024646 
+ SKY130_FD_PR__ESD_NFET_01V8__VSAT_DIFF_0=29832.0 SKY130_FD_PR__ESD_NFET_01V8__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__NFACTOR_DIFF_0=0.3284 SKY130_FD_PR__ESD_NFET_01V8__B1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__UA_DIFF_1=1.1282e-10 
+ SKY130_FD_PR__ESD_NFET_01V8__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITSD_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__TVOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__VOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__K2_DIFF_1=-0.017137 
+ SKY130_FD_PR__ESD_NFET_01V8__UB_DIFF_1=2.3412e-19 SKY130_FD_PR__ESD_NFET_01V8__VTH0_DIFF_1=0.055271 
+ SKY130_FD_PR__ESD_NFET_01V8__U0_DIFF_1=0.0037507 SKY130_FD_PR__ESD_NFET_01V8__VSAT_DIFF_1=15696.0 
+ SKY130_FD_PR__ESD_NFET_01V8__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__NFACTOR_DIFF_1=-0.27022 
+ SKY130_FD_PR__ESD_NFET_01V8__B1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__B0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__B0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__AGS_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__UA_DIFF_2=1.2882e-10 SKY130_FD_PR__ESD_NFET_01V8__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITS_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PCLM_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__K2_DIFF_2=-0.0077745 SKY130_FD_PR__ESD_NFET_01V8__UB_DIFF_2=-2.6082e-19 
+ SKY130_FD_PR__ESD_NFET_01V8__VTH0_DIFF_2=0.056219 SKY130_FD_PR__ESD_NFET_01V8__U0_DIFF_2=0.0018148 
+ SKY130_FD_PR__ESD_NFET_01V8__VSAT_DIFF_2=26605.0 SKY130_FD_PR__ESD_NFET_01V8__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__NFACTOR_DIFF_2=-0.44799 SKY130_FD_PR__ESD_NFET_01V8__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__RDSW_DIFF_2=0.0
*
* sky130_fd_pr__esd_nfet_01v8, Bin 000, W = 20.35, L = 0.165
* ----------------------------------------
*
* sky130_fd_pr__esd_nfet_01v8, Bin 001, W = 40.31, L = 0.165
* ----------------------------------------
*














* sky130_fd_pr__esd_nfet_01v8, Bin 002, W = 5.4, L = 0.18
* -------------------------------------
.INCLUDE sky130_fd_pr__esd_nfet_01v8.pm3.spice




















