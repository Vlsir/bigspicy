** Translated using xdm 2.6.0 on Nov_14_2022_16_05_13_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_B__TOXE_MULT=1.0365 SKY130_FD_PR__RF_NFET_01V8_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_NFET_01V8_B__OVERLAP_MULT=0.98 SKY130_FD_PR__RF_NFET_01V8_B__AJUNCTION_MULT=1.1505 
+ SKY130_FD_PR__RF_NFET_01V8_B__PJUNCTION_MULT=1.1793 SKY130_FD_PR__RF_NFET_01V8_B__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__RF_NFET_01V8_B__WINT_DIFF=2.252e-8 SKY130_FD_PR__RF_NFET_01V8_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__DLC_DIFF=-11.107e-9 SKY130_FD_PR__RF_NFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__XGW_DIFF=4.504e-8 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_0=0.016061 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_0=7256.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_0=0.0079631 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_0=-0.0019138 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_1=0.020817 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_1=9830.4 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_1=0.014994 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_1=-0.002237 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_2=0.0086842 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_2=19450.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_2=0.032627 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_2=-0.0030221 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_3=0.025003 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_3=1653.2 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_3=0.0026575 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_3=-0.0083307 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_4=0.00020419 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_4=12334.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_4=0.015143 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_4=-0.0053582 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_5=0.0016884 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_5=11246.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_5=0.034079 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_5=-0.0028787 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_6=-0.006203 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_6=0.0065467 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_6=-4610.9 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_6=0.001022 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_7=0.013198 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_7=-0.0055047 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_7=-0.0028156 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_7=9383.7 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_8=0.031946 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_8=-0.0050561 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_8=-0.0043506 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_8=12165.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_0=0.0068964 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_0=-0.0035814 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_0=0.040659 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_0=-2843.6 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_1=0.019365 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_1=-0.0039029 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_1=0.0080414 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_1=11376.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_2=0.035011 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_2=-0.0035828 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_2=0.0072093 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_2=24875.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_3=526.28 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_3=0.0028165 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_3=-0.0086312 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_3=0.018526 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_4=14947.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_4=0.017688 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_4=-0.008178 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_4=-0.0046622 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_5=40210.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_5=0.035635 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_5=-0.0070625 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_5=-0.0049699 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_6=-4885.3 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_6=0.0013795 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_6=-0.0060867 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_6=0.0069395 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_7=-0.0068351 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_7=3065.3 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_7=0.016371 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_7=-0.012469 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_8=-0.0078852 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_8=-0.0064297 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_8=34241.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_8=0.033541
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*





* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_b.pm3.spice














