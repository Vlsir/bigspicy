** Translated using xdm 2.6.0 on Nov_14_2022_16_05_33_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 9
.PARAM 
+ SKY130_FD_PR__NFET_03V3_NVT__TOXE_MULT=1.0 SKY130_FD_PR__NFET_03V3_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_03V3_NVT__OVERLAP_MULT=0.77117 SKY130_FD_PR__NFET_03V3_NVT__AJUNCTION_MULT=0.97602 
+ SKY130_FD_PR__NFET_03V3_NVT__PJUNCTION_MULT=1.0437 SKY130_FD_PR__NFET_03V3_NVT__LINT_DIFF=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__WINT_DIFF=0.0 SKY130_FD_PR__NFET_03V3_NVT__DLC_DIFF=-1.5781e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__DWC_DIFF=0.0 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_0=0.038449 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_0=0.0019135 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_0=-1.3838 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_0=-0.015836 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_0=-0.00065697 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_0=-3837.2 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_0=-1.4132e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_0=3.4977e-11 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_1=5.3407e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_1=0.033082 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_1=0.0096743 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_1=-1.3958 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_1=-0.015324 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_1=-0.0011594 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_1=-6763.8 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_1=1.0429e-19 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_2=2.6095e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_2=5.8204e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_2=0.0057767 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_2=-0.46503 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_2=0.0032323 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_2=0.0063254 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_2=-4056.8 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_3=-3.3361e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_3=3.7397e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_3=0.040673 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_3=0.0032721 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_3=-1.3621 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_3=-0.01875 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_3=-0.00011074 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_3=-4396.2 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_4=3.7224e-19 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_4=2.2268e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_4=0.045453 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_4=0.010004 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_4=-1.3404 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_4=-0.018338 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_4=-0.0018856 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_4=-8376.1 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_5=0.011241 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_5=-6843.2 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_5=3.0597e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_5=7.2969e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_5=0.012715 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_5=-1.6434 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_5=0.051876 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_6=-0.746 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_6=0.022008 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_6=0.007881 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_6=-3534.9 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_6=2.3973e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_6=8.5737e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_6=0.012066 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_7=0.04193 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_7=0.011117 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_7=-1.3436 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_7=-0.014154 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_7=-0.0017689 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_7=-7893.2 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_7=2.6547e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_7=4.0061e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_8=0.0084797 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_8=-0.43724 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_8=-0.0034771 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_8=0.005952 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_8=-5528.9 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_8=2.4645e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_8=5.5525e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_8=0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
*














* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_03v3_nvt.pm3.spice




















