** Translated using xdm 2.6.0 on Nov_14_2022_16_05_16_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__RF_PFET_01V8_B__TOXE_MULT=0.948 SKY130_FD_PR__RF_PFET_01V8_B__RBPB_MULT=0.8 
+ SKY130_FD_PR__RF_PFET_01V8_B__OVERLAP_MULT=0.95436 SKY130_FD_PR__RF_PFET_01V8_B__AJUNCTION_MULT=0.90161 
+ SKY130_FD_PR__RF_PFET_01V8_B__PJUNCTION_MULT=0.90587 SKY130_FD_PR__RF_PFET_01V8_B__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__RF_PFET_01V8_B__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__RF_PFET_01V8_B__RSHG_DIFF=-7.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__DLC_DIFF=1.7325e-8 SKY130_FD_PR__RF_PFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__XGW_DIFF=-6.4250e-8 SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT=0.85 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT=0.77 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT=0.77 
+ SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT_2=0.85 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT_2=0.80 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT_2=0.80 SKY130_FD_PR__RF_PFET_01V8__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RS_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_0=0.0036576 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_0=-0.00034614 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_0=-0.092407 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_0=-19636.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_1=-0.0076806 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_1=-0.00019683 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_1=-0.079373 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_1=-15546.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_2=-0.033345 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_2=-3.0791e-5 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_2=-0.030098 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_2=-6434.1 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_3=-0.0012925 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_3=-0.00028011 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_3=-0.12131 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_3=-18686.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_4=0.00024736 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_4=-0.00041476 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_4=-0.071611 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_4=-11333.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_5=-0.016582 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_5=-0.00016695 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_5=-0.025831 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_5=-1107.2 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_6=-0.0014721 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_6=-0.00053506 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_6=-0.13112 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_6=-16484.0 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_7=-0.00025473 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_7=-17993.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_7=0.00033491 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_7=-0.077674 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_8=-0.035077 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_8=-0.00020922 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_8=-5719.7 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_8=-0.019564 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_0=0.0065905 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_0=-0.00050702 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_0=-0.081008 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_0=-20196.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_1=-0.0063812 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_1=-0.00027314 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_1=-0.065695 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_1=-12293.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_2=-7.2735e-5 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_2=-0.022778 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_2=272.66 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_2=-0.034415 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_3=0.00078898 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_3=-0.0003818 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_3=-0.11908 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_3=-16139.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_4=-0.00058216 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_4=-0.058416 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_4=-11485.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_4=0.0039762 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_5=-0.01803 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_5=-0.00025609 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_5=-7303.4 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_5=-0.016473 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_6=-0.12568 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_6=-0.00035343 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_6=-16543.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_6=0.00030278 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_7=0.0028314 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_7=-0.073523 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_7=-0.000511 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_7=-15224.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_8=-0.018202 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_8=-0.022497 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_8=-0.00030626 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_8=4136.5 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_8=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_pfet_01v8_b.pm3.spice














