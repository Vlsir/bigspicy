** Translated using xdm 2.6.0 on Nov_14_2022_16_05_35_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
* Number of bins: 1
.PARAM 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__TOX_MULT=1.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__AJUNCTION_MULT=9.9543e-1 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__PJUNCTION_MULT=1.0204e+0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__OVERLAP_MULT=0.89805 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__LINT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__WINT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DWG_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__K3_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DVT0_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DVT0W_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__NLX_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CIT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CDSC_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CDSCB_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CDSCD_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT2_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT1L_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DLC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DWC_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__K2_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__U0_DIFF_0=0.0027584 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VSAT_DIFF_0=3855.4 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VTH0_DIFF_0=-0.15663 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT1_DIFF_1=3.8227e-2 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__NFACTOR_DIFF_1=1.4138e-1 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VOFF_DIFF_1=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__K2_DIFF_1=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__U0_DIFF_1=1.2956e-3 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VSAT_DIFF_1=1.3679e+4 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VTH0_DIFF_1=-5.7093e-3
*


* sky130_fd_pr__special_nfet_pass_flash, Bin 000, W = 0.45, L = 0.15
* -----------------------------------
*







* sky130_fd_pr__special_nfet_pass_flash, Bin 001, W = 0.35, L = 0.15
* -----------------------------------
* Number of bins: 1







.PARAM 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__TOX_MULT=1.0 SKY130_FD_PR__SPECIAL_NFET_PASS__AJUNCTION_MULT=9.9543e-1 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__PJUNCTION_MULT=1.0204e+0 SKY130_FD_PR__SPECIAL_NFET_PASS__OVERLAP_MULT=0.9842 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__LINT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__WINT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__K3_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__DVT0_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__CIT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__CDSC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__CDSCB_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__CDSCD_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__KT2_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__KT1L_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__DLC_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__DWC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__KT1_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__VSAT_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__K2_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__U0_DIFF_0=-0.0029226 SKY130_FD_PR__SPECIAL_NFET_PASS__VTH0_DIFF_0=0.027522 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__RDSW_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__VOFF_DIFF_0=0.0
*




* sky130_fd_pr__special_nfet_pass, Bin 000, W = 0.14, L = 0.15
* ----------------------------------
* Number of bins: 1








.PARAM 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__TOX_MULT=1.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__AJUNCTION_MULT=9.9543e-1 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__PJUNCTION_MULT=1.0204e+0 SKY130_FD_PR__SPECIAL_NFET_LATCH__OVERLAP_MULT=0.9842 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__LINT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__WINT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__K3_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__DVT0_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__DVT1_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__CIT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__CDSC_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__CDSCB_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__CDSCD_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__KT2_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__DLC_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__DWC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__VOFF_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__RDSW_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__K2_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__U0_DIFF_0=0.00030368 SKY130_FD_PR__SPECIAL_NFET_LATCH__VTH0_DIFF_0=0.020952 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__VSAT_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__NFACTOR_DIFF_0=0.0
*




* sky130_fd_pr__special_nfet_latch, Bin 000, W = 0.21, L = 0.15
* --------------------------------
* Number of bins: 1








.PARAM 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__TOX_MULT=1.0 SKY130_FD_PR__SPECIAL_PFET_PASS__AJUNCTION_MULT=9.9626e-1 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__PJUNCTION_MULT=1.0009e+0 SKY130_FD_PR__SPECIAL_PFET_PASS__OVERLAP_MULT=9.5435e-1 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__LINT_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__WINT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__K3_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__DVT0_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__CIT_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__CDSC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__CDSCB_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__CDSCD_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__KT2_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__KT1L_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__DLC_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__DWC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__VOFF_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__VSAT_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__VTH0_DIFF_0=0.0081943 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__K2_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__U0_DIFF_0=-0.00044468 SKY130_FD_PR__SPECIAL_PFET_PASS__RDSW_DIFF_0=0.0
*




* sky130_fd_pr__special_pfet_pass, Bin 000, W = 0.14, L = 0.15
* --------------------------------
.INCLUDE sky130_fd_pr__special_nfet_latch__mismatch.corner.spice








.INCLUDE sky130_fd_pr__special_nfet_pass__mismatch.corner.spice
.INCLUDE sky130_fd_pr__special_nfet_pass_flash__mismatch.corner.spice
.INCLUDE sky130_fd_pr__special_pfet_pass__mismatch.corner.spice
.INCLUDE sky130_fd_pr__special_nfet_pass_lvt__tt.corner.spice
