** Translated using xdm 2.6.0 on Nov_14_2022_16_05_35_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TOXE_MULT=1.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RSHN_MULT=1.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__OVERLAP_MULT=0.89805 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AJUNCTION_MULT=9.9505e-1 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PJUNCTION_MULT=1.0144e+0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__LINT_DIFF=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__WINT_DIFF=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__DLC_DIFF=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__DWC_DIFF=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_0=0.23362 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_0=0.010406 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_0=0.001245 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_0=0.012769 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_0=-1672.2 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_0=2.4153e-19 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_0=-8.8395e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_1=0.23014 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_1=0.010327 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_1=0.0029959 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_1=0.014049 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_1=-1443.7 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_1=3.4221e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_1=-2.42e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_2=0.23391 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_2=0.010304 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_2=0.0012741 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_2=0.013326 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_2=-43.451 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_2=3.291e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_2=-7.333e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_3=-1.7201e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_3=0.23086 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_3=0.010034 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_3=0.0010628 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_3=0.01319 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_3=33.54 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_3=3.183e-19 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_4=2.7249e-19 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_4=-7.6527e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_4=0.22609 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_4=0.0099796 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_4=0.0013927 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_4=0.011469 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_4=-907.07 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_5=-6.1783e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_5=8.2128e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_5=0.27056 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_5=-0.021325 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_5=-0.26694 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_5=0.047533 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_5=-0.0063931 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_5=0.010431 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_6=6.0666e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_6=-7.0128e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_6=0.22669 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_6=0.010019 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_6=0.0016874 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_6=0.011396 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_6=1500.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_7=3019.2 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_7=9.7977e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_7=3.2228e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_7=0.19932 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_7=0.010207 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_7=0.0014468 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_7=0.011899 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_8=-0.0088519 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_8=-8.0124e-5 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_8=-6.7671e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_8=5.5348e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_8=0.25888 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_8=0.0071088 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_8=0.0024548 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_8=0.010977 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_9=0.0014488 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_9=0.0037985 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_9=0.002943 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_9=-191.5 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_9=1.3051e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_9=-1.3283e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_9=0.20721 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_10=2.8803e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_10=-2502.2 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_10=8.2506e-20 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_10=0.0031768 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_10=0.29591 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_10=-0.00045045 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_10=0.013543 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
*
















* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
.INCLUDE sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice























