** Translated using xdm 2.6.0 on Nov_14_2022_16_05_35_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_MULT=1.0 SKY130_FD_PR__NFET_05V0_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_05V0_NVT__OVERLAP_MULT=7.7117e-1 SKY130_FD_PR__NFET_05V0_NVT__AJUNCTION_MULT=9.7602e-1 
+ SKY130_FD_PR__NFET_05V0_NVT__PJUNCTION_MULT=1.0437e+0 SKY130_FD_PR__NFET_05V0_NVT__LINT_DIFF=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__WINT_DIFF=0.0 SKY130_FD_PR__NFET_05V0_NVT__DLC_DIFF=-1.5781e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__DWC_DIFF=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_0=0.010308 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_0=0.0064317 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_0=-0.00025708 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_0=-0.0078378 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_0=-2.691e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_0=-0.0046033 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_0=0.00034013 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_0=-1.3689e-18 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_1=-1.2472e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_1=0.029952 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_1=-0.00044213 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_1=-0.0039719 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_1=-0.0070434 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_1=-2.4351e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_1=-0.0022002 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_1=-0.00056708 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_2=-1.5224e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_2=-0.044586 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_2=0.0015915 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_2=-0.008363 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_2=-3.3419e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_2=-2848.5 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_2=-0.0011931 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_3=-1.6915e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_3=0.0075894 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_3=-9.6861e-19 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_3=0.064023 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_3=0.0012767 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_3=-0.0046305 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_3=-0.0066322 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_3=-0.013446 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_4=-0.0078468 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_4=-0.0057166 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_4=-2.429e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_4=-0.0084686 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_4=-1.2894e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_4=0.024393 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_4=-0.035687 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_4=-0.0016893 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_5=-0.00013553 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_5=-0.0079399 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_5=-0.0050535 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_5=-2.1501e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_5=0.0053237 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_5=-1.2037e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_5=0.053081 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_5=0.02762 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_6=0.00043703 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_6=-0.0023615 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_6=-0.0068188 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_6=-0.011078 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_6=-1.9014e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_6=-0.00041719 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_6=-1.0585e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_6=0.055346 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_7=0.0016268 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_7=0.00035232 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_7=-0.0094947 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_7=-0.014254 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_7=-2.898e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_7=-3146.5 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_7=-1.429e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_8=0.017467 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_8=8.0096e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_8=-0.0049283 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_8=-0.0086023 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_8=-0.031553 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_8=-2.2873e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_8=1.6514e-9 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_8=-1.2296e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_9=-0.011611 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_9=-0.0030036 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_9=-0.0089225 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_9=-0.010333 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_9=-1.3766e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_9=-6052.7 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_9=-9.127e-19 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_10=-4889.9 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_10=-0.010495 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_10=0.011275 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_10=-0.0096426 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_10=0.00063457 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_10=-2.505e-11 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_10=-1.3111e-18 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0, L = 2.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0, L = 4.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0, L = 0.9
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0, L = 25.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0, L = 2.0
* ------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0, L = 4.0
* ------------------------------------
*














* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0, L = 8.0
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0, L = 0.9
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42, L = 1.0
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42, L = 0.9
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7, L = 0.9
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_05v0_nvt.pm3.spice




















