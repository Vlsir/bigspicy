** Translated using xdm 2.6.0 on Nov_14_2022_16_05_34_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__RF_PFET_01V8_B__TOXE_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_B__RBPB_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__OVERLAP_MULT=9.5435e-1 SKY130_FD_PR__RF_PFET_01V8_B__AJUNCTION_MULT=9.9626e-1 
+ SKY130_FD_PR__RF_PFET_01V8_B__PJUNCTION_MULT=1.0009 SKY130_FD_PR__RF_PFET_01V8_B__LINT_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__WINT_DIFF=0.0 SKY130_FD_PR__RF_PFET_01V8_B__RSHG_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__DLC_DIFF=0.0 SKY130_FD_PR__RF_PFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__XGW_DIFF=0.0 SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT_2=1.0 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT_2=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT_2=1.0 SKY130_FD_PR__RF_PFET_01V8__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RS_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_0=-0.023953 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_0=-0.00025608 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_0=0.0054151 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_0=-1792.7 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_1=-0.0146 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_1=-0.00017534 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_1=-0.0013289 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_1=-3939.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_2=-0.017504 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_2=-0.00011528 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_2=0.0016874 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_2=-3705.2 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_3=-0.025672 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_3=-0.00043953 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_3=0.00554 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_3=-7604.3 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_4=-0.016429 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_4=-0.00040298 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_4=0.0090164 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_4=222.9 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_5=-0.018578 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_5=-0.00022966 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_5=0.0043185 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_5=12358.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_6=-0.026387 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_6=-0.00078906 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_6=0.013291 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_6=-3996.4 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_7=-0.00030611 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_7=-5407.7 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_7=-0.013695 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_7=0.0054619 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_8=0.0030552 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_8=-0.00032694 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_8=2232.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_8=-0.017831 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_0=-0.022271 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_0=-0.00043404 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_0=0.018047 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_0=-1656.1 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_1=-0.014049 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_1=-0.0002533 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_1=0.012426 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_1=876.35 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_2=-0.0001857 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_2=0.0094773 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_2=15921.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_2=-0.018595 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_3=-0.023461 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_3=-0.00053503 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_3=0.0064872 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_3=-2980.8 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_4=-0.00062465 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_4=0.022342 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_4=-1155.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_4=-0.012789 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_5=0.012097 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_5=-0.00033445 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_5=9117.5 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_5=-0.018599 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_6=0.017753 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_6=-0.00064602 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_6=-2850.2 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_6=-0.0251 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_7=-0.010953 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_7=0.0097164 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_7=-0.00057548 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_7=-3914.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_8=-0.016606 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_8=0.015491 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_8=-0.00044041 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_8=11410.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_8=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_pfet_01v8_b.pm3.spice














