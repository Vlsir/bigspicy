** Translated using xdm 2.6.0 on Nov_14_2022_16_05_29_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10 w = 3.01 l = 0.50 m = 10 ad = 0.421 pd = 3.29 as = 0.51 ps = 3.948 nrd = 40.44 nrs = 33.70 mult = {10*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10 w = 3.01 l = 0.50 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04 w = 3.01 l = 0.50 m = 4 ad = 0.421 pd = 3.29 as = 0.63 ps = 4.935 nrd = 40.44 nrs = 26.96 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04 w = 3.01 l = 0.50 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00 l = 0.50 m = 10 ad = 0.707 pd = 5.33 as = 0.85 ps = 6.396 nrd = 24.27 nrs = 20.22 mult = {10*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00 l = 0.50 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00 l = 0.50 m = 4 ad = 0.707 pd = 5.33 as = 1.06 ps = 7.995 nrd = 24.267 nrs = 16.178 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00 l = 0.50 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00 l = 0.50 m = 10 ad = 0.993 pd = 7.37 as = 1.19 ps = 8.844 nrd = 17.33 nrs = 14.44 mult = {10*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00 l = 0.50 m = 2 ad = 2.127 pd = 14.78 as = 0.0 ps = 0.0 nrd = 8.67 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00 l = 0.50 m = 4 ad = 0.993 pd = 7.37 as = 1.49 ps = 11.055 nrd = 17.33 nrs = 11.56 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00 l = 0.50 m = 2 ad = 2.127 pd = 14.78 as = 0.0 ps = 0.0 nrd = 8.67 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00 l = 0.50 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 24.267 nrs = 12.133 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00 l = 0.50 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50
.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM02 w = 3.01 l = 0.50 m = 2 ad = 0.42 pd = 3.29 as = 0.84 ps = 6.58 nrd = 40.44 nrs = 20.22 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50_dummy b b s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM02 w = 3.01 l = 0.50 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50
