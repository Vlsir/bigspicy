** Translated using xdm 2.6.0 on Nov_14_2022_16_05_04_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

*.param
* .model sky130_fd_pr__nfet_20v0_nvt__parasitic__diode_ps2dn d  level = 3.0   tlevc = 1.0   scalm = 1.0e-6   area = 1.0e+12   cj = '1.6920e-004*sky130_fd_pr__nfet_20v0__cjdnwpsubjunction_mult*1e-12*sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult' ; Units: farad/meter^2   mj = '0.56056*sky130_fd_pr__nfet_20v0__mjdnwpsubjunction_mult'   pb = '0.21294*sky130_fd_pr__nfet_20v0__pbdnwpsubjunction_mult' ; Units: volt   cjsw = '8.1380e-010*sky130_fd_pr__nfet_20v0__cjdnwpsubjunction_mult*1e-6*sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult' ; Units: farad/meter   mjsw = '0.18742*sky130_fd_pr__nfet_20v0__mjdnwpsubjunction_mult'   php = '0.21294*sky130_fd_pr__nfet_20v0__pbdnwpsubjunction_mult' ; Units: volt   cta = 0.0031223 ; Units: 1/coulomb   ctp = 0.0014703 ; Units: 1/coulomb   tpb = 0.0016859 ; Units: volt/coulomb   tphp = 0.0016859 ; Units: volt/coulomb   js = 6.1049e-017 ; Units: amper/meter^2   jsw = 8.1115e-016 ; Units: amper/meter   n = 1.0791   rs = 900 ; Units: ohm (ohm/meter^2 if area defined)   ik = '2.08e-009/1e-12' ; Units: amper/meter^2   ikr = '0/1e-12' ; Units: amper/meter^2   vb = 'sky130_fd_pr__nfet_20v0__vb' ; Units: volt   ibv = 0.00106 ; Units: amper   trs = 0 ; Units: 1/coulomb   eg = 1.17 ; Units: electron-volt   xti = 1.0   tref = 30 ; Units: coulomb   tcv = 0 ; Units: 1/coulomb   gap1 = 0.000473 ; Units: electron-volt/coulomb   gap2 = 1110.0   ttt1 = 0 ; Units: 1/coulomb   ttt2 = 0 ; Units: 1/coulomb^2   tm1 = 0 ; Units: 1/coulomb   tm2 = 0 ; Units: 1/coulomb^2   lm = 0 ; Units: meter   lp = 0 ; Units: meter   wm = 0 ; Units: meter   wp = 0 ; Units: meter   xm = 0 ; Units: meter   xoi = 10000.0   xom = 10000 ; Units: angstrom   xp = 0 ; Units: meter   xw = 0 ; Units: meter; HSpice Parser Retained (as a comment). Continuing.
* Junction Capacitance Parameters




* Diode IV Parameters










* Default Parameters












