** Translated using xdm 2.6.0 on Nov_14_2022_16_05_18_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_MULT=0.9635 SKY130_FD_PR__NFET_05V0_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_05V0_NVT__OVERLAP_MULT=5.1025e-1 SKY130_FD_PR__NFET_05V0_NVT__AJUNCTION_MULT=6.8772e-1 
+ SKY130_FD_PR__NFET_05V0_NVT__PJUNCTION_MULT=9.0190e-1 SKY130_FD_PR__NFET_05V0_NVT__LINT_DIFF=1.21275e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__WINT_DIFF=-2.252e-8 SKY130_FD_PR__NFET_05V0_NVT__DLC_DIFF=1.6112e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__DWC_DIFF=-2.252e-8 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_0=0.056665 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_0=-0.052927 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_0=-0.00059672 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_0=-0.0090633 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_0=-3.141e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_0=-0.030851 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_0=-0.005637 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_0=-1.5907e-18 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_1=-1.357e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_1=-0.019967 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_1=-0.032965 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_1=-0.0051327 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_1=-0.0077525 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_1=-2.636e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_1=-0.018137 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_1=-0.0051202 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_2=-1.8782e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_2=0.066292 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_2=0.00087158 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_2=-0.0096682 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_2=-4.2384e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_2=-6160.2 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_2=-0.03046 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_3=-2.0373e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_3=-0.0020789 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_3=-1.0928e-18 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_3=0.015653 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_3=0.0012297 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_3=-0.0052343 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_3=-0.0065532 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_3=-0.024011 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_4=-0.0083037 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_4=-0.020154 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_4=-2.6021e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_4=-0.038115 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_4=-1.4421e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_4=-0.05753 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_4=-0.17718 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_4=-0.0022264 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_5=-0.00093844 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_5=-0.007664 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_5=-0.017363 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_5=-2.4895e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_5=-0.0093971 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_5=-1.3242e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_5=-0.0035696 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_5=-0.044469 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_6=-0.047321 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_6=-0.0028201 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_6=-0.0068477 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_6=-0.023509 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_6=-2.2313e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_6=-0.009358 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_6=-1.1832e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_6=-0.022424 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_7=0.043963 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_7=-3.5325e-6 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_7=-0.010425 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_7=-0.038579 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_7=-3.6456e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_7=-6428.9 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_7=-1.7165e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_8=0.017354 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_8=1.5203e-7 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_8=-0.0095342 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_8=-0.0085304 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_8=-0.055166 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_8=-3.4036e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_8=-4.5502e-9 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_8=-1.6434e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_9=-0.13265 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_9=-0.0070168 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_9=-0.0087887 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_9=-0.042098 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_9=-2.2834e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_9=-8459.3 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_9=-1.3613e-18 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_10=-7916.1 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_10=-0.035797 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_10=0.028686 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_10=-0.010001 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_10=0.00041829 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_10=-3.5554e-11 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_10=-1.6633e-18 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0, L = 2.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0, L = 4.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0, L = 0.9
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0, L = 25.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0, L = 2.0
* ------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0, L = 4.0
* ------------------------------------
*














* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0, L = 8.0
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0, L = 0.9
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42, L = 1.0
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42, L = 0.9
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7, L = 0.9
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_05v0_nvt.pm3.spice




















