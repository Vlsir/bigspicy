** Translated using xdm 2.6.0 on Nov_14_2022_16_05_08_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__cap_mim_m3_1 c0 c1 PARAMS: W=1 L=1 MF=1
.PARAM WC='w+m3_dw*1e6+tol_m3*1e6'
.PARAM LC='l+m3_dw*1e6+tol_m3*1e6'
.PARAM VIA3_SPACING='(0.17+0.25+0.140)*(0.17+0.25+0.140)'
.PARAM NUM_CONTACTS='(wc*lc/via3_spacing)'
.PARAM R1='rm3*(lc)/(wc)'
.PARAM R2='rcvia3/num_contacts'
.PARAM CAREA='camimc*(wc)*(lc)'
.PARAM CPERIM='cpmimc*((wc)+(lc))*2'
.PARAM 
+ CZERO='carea + cperim+MC_MM_SWITCH*AGAUSS(0,1.0,1)*0.01*2.8*(carea + cperim)/sqrt(wc*lc*mf)'
C1 c0 a TC1=0 TC2=0.0 C='czero'
* rs1 a        b1 'r1' tc1 = {tc1rm3} tc2 = {tc2rm3}; HSpice Parser Retained (as a comment). Continuing.
* rs2 b1        c1 'r2' tc1 = {tc1rvia3} tc2 = {tc2rvia3}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__cap_mim_m3_1
