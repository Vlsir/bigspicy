** Translated using xdm 2.6.0 on Nov_14_2022_16_05_29_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
.PARAM 
+ CAPUNITS=1.0e-6 DKISEPP5X=0.745 DKNFPP=1.0 DKNFPP5X=1.0009 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CDSC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CDSCB_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CDSCD_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__CIT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DVT0_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DVT0W_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__DWG_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__K2_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__K2_DIFF_1=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__K3_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT1_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT1L_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__KT2_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__LINT_SLOPE=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__NFACTOR_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__NLX_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__TOX_SLOPE=0.006589 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VOFF_SLOPE=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__VTH0_SLOPE=0.010889 SKY130_FD_PR__SPECIAL_NFET_PASS_FLASH__WINT_SLOPE=0.0 
+ GLOBALK=1.0 HV_DLC_ROTWEAK=0.0 LOCALKSWITCH=1.0 LV_DLC_ROTWEAK=0.0 LVHVT_DLC_ROTWEAK=0.0 
+ LVT_DLC_ROTWEAK=0.0 MCL1P1F_CC_W_1_200_S_5_250=0.0 MCM1L1D_CC_W_1_360_S_0_360=3.25e-11 
+ MCM2D_CC_W_0_140_S_1_540=2.6e-11 MCM2M1L1_CC_W_1_120_S_3_500=5.0e-14 MCM2P1F_CC_W_1_200_S_0_420=4.11e-11 
+ MCM3M2_CC_W_0_300_S_3_300=9.9e-12 MCM4M2F_CF_W_1_120_S_0_140=2.69e-12 MCM5M1P1_CC_W_0_140_S_0_840=3.22e-11 
+ MCM5M2F_CC_W_1_120_S_0_840=4.63e-11 MCM5M4_CC_W_1_600_S_10_000=4.0e-12 MCM5M4M3_CC_W_2_400_S_9_000=5.0e-14 
+ MCRDLM3M2_CC_W_0_300_S_2_100=1.55e-11 MCRDLM4L1_CC_W_0_300_S_3_300=1.91e-11 MCRDLM4P1_CC_W_0_300_S_3_300=2.02e-11 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_44=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGIDL_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_22=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_24=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_8=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_22=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_24=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_44=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_8=0.0 SKY130_FD_PR__NFET_G5V0D10V5__BGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__ETA0_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_22=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_24=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_44=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_8=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KETA_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__KU0_DIFF=-4.5e-8 
+ SKY130_FD_PR__NFET_G5V0D10V5__KVSAT_DIFF=0.3 SKY130_FD_PR__NFET_G5V0D10V5__KVTH0_DIFF=1.1e-8 
+ SKY130_FD_PR__NFET_G5V0D10V5__LINT_SLOPE=0.0 SKY130_FD_PR__NFET_G5V0D10V5__LKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__LKVTH0_DIFF=0.0 SKY130_FD_PR__NFET_G5V0D10V5__NFACTOR_SLOPE=0.12 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PCLM_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_22=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_24=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_44=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__PDITSD_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_22=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_24=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_44=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_G5V0D10V5__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__B_LINT_SLOPE=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5__B_NFACTOR_SLOPE=0.12 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__B_TOXE_SLOPE=0.008 SKY130_FD_PR__RF_NFET_G5V0D10V5__B_TOXE_SLOPE1=0.0205 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__B_TOXE_SLOPE2=0.01 SKY130_FD_PR__RF_NFET_G5V0D10V5__B_TOXE_SLOPE3=0.0067 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__B_VOFF_SLOPE=0.13 SKY130_FD_PR__RF_NFET_G5V0D10V5__B_VTH0_SLOPE=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__B_WINT_SLOPE=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__BASE__DLC_ROTWEAK=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__PCLM_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5__LINT1_SLOPE=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__LINT_SLOPE=3.0e-9 SKY130_FD_PR__RF_NFET_G5V0D10V5__NFACTOR_SLOPE=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX2_SLOPE=0.0086 SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX3_SLOPE=0.0055 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX4_SLOPE=0.0255 SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX_OFFSET=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX_SLOPE=0.008 SKY130_FD_PR__RF_NFET_G5V0D10V5__VOFF2_SLOPE=0.0085 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5__VOFF_SLOPE=0.00375 SKY130_FD_PR__RF_NFET_G5V0D10V5__WINT_SLOPE=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__RSHN_MULT=1.0 SKY130_FD_PR__NFET_G5V0D10V5__TOXE_SLOPE=0.008 
+ SKY130_FD_PR__NFET_G5V0D10V5__TOXE_SLOPE1=0.0205 SKY130_FD_PR__NFET_G5V0D10V5__TOXE_SLOPE2=0.01 
+ SKY130_FD_PR__NFET_G5V0D10V5__TOXE_SLOPE3=0.0067 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_11=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_13=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_15=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_20=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_22=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_24=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_26=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_28=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_33=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_40=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_42=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_44=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_46=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_48=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_G5V0D10V5__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_12=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_16=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_18=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_21=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_27=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_29=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_30=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_32=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_34=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_36=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_38=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_41=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_47=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VOFF_SLOPE=0.13 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_14=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_17=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_19=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_23=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_25=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_31=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_35=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_37=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_39=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_43=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_45=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_7=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__VSAT_DIFF_9=0.0 SKY130_FD_PR__NFET_G5V0D10V5__VTH0_SLOPE=0.0 
+ SKY130_FD_PR__NFET_G5V0D10V5__WINT_SLOPE=0.0 SKY130_FD_PR__NFET_G5V0D10V5__WKU0_DIFF=2.0e-7 
+ SKY130_FD_PR__NFET_G5V0D10V5__WKVTH0_DIFF=6.5e-7 SKY130_FD_PR__NFET_G5V0D10V5__WLOD_DIFF=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RSHN_MULT=1.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__DLC_ROTWEAK={hv_dlc_rotweak} SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KU0_DIFF=-3.0e-8 SKY130_FD_PR__NFET_05V0_NVT__KVSAT_DIFF=0.4 
+ SKY130_FD_PR__NFET_05V0_NVT__KVTH0_DIFF=-7.0e-9 SKY130_FD_PR__NFET_05V0_NVT__LINT_SLOPE=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__LKU0_DIFF=0.0 SKY130_FD_PR__NFET_05V0_NVT__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_SLOPE=0.02 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_SLOPE=0.00105 SKY130_FD_PR__NFET_05V0_NVT__TOXE_SLOPE1=0.01205 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_SLOPE2=0.02525 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_SLOPE=0.0035 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_SLOPE=0.0012 
+ SKY130_FD_PR__NFET_05V0_NVT__WINT_SLOPE=0.0 SKY130_FD_PR__NFET_05V0_NVT__WKU0_DIFF=2.0e-7 
+ SKY130_FD_PR__NFET_05V0_NVT__WKVTH0_DIFF=8.0e-7 SKY130_FD_PR__NFET_05V0_NVT__WLOD_DIFF=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B0_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8_LVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__DLC_ROTWEAK={lvt_dlc_rotweak} SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__ETA0_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__KU0_DIFF=-2.7e-8 
+ SKY130_FD_PR__NFET_01V8_LVT__KVSAT_DIFF=0.2 SKY130_FD_PR__NFET_01V8_LVT__KVTH0_DIFF=7.9e-9 
+ SKY130_FD_PR__NFET_01V8_LVT__LINT_SLOPE=0.0 SKY130_FD_PR__NFET_01V8_LVT__LKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__LKVTH0_DIFF=0.0 SKY130_FD_PR__NFET_01V8_LVT__NFACTOR_SLOPE=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8_LVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8_LVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8_LVT__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RD_MULT=1.0 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RS_MULT=1.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__B_TOXE_SLOPE=0.003443 SKY130_FD_PR__RF_NFET_01V8_LVT__B_VTH0_SLOPE=0.006056 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__DWC_DIFF=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT__BASE__DLC_ROTWEAK=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__TOXE1_SLOPE=0.008089 SKY130_FD_PR__RF_NFET_01V8_LVT__TOXE_SLOPE=0.006789 
+ SKY130_FD_PR__NFET_01V8_LVT__RSHN_MULT=1.0 SKY130_FD_PR__NFET_01V8_LVT__TOXE_SLOPE=0.003443 
+ SKY130_FD_PR__NFET_01V8_LVT__TOXE_SLOPE1=0.002443 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__VOFF_SLOPE=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__VSAT_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8_LVT__VTH0_SLOPE=0.005456 
+ SKY130_FD_PR__NFET_01V8_LVT__VTH0_SLOPE1=0.005456 SKY130_FD_PR__NFET_01V8_LVT__VTH0_SLOPE2=0.007456 
+ SKY130_FD_PR__NFET_01V8_LVT__WINT_SLOPE=0.0 SKY130_FD_PR__NFET_01V8_LVT__WKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_01V8_LVT__WKVTH0_DIFF=3.0e-7 SKY130_FD_PR__NFET_01V8_LVT__WLOD_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__K2_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__UA_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__UB_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__VOFF_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__CDSC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__CDSCB_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__CDSCD_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__CIT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__DLC_ROTWEAK={lv_dlc_rotweak} 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__DVT0_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__K2_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__K3_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__KT1L_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__KT2_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__LINT_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__NFACTOR_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__TOX_SLOPE=0.003589 SKY130_FD_PR__SPECIAL_NFET_PASS__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__VOFF_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS__VTH0_SLOPE=0.005589 SKY130_FD_PR__SPECIAL_NFET_PASS__WINT_SLOPE=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LOWLEAKAGE__DLC_ROTWEAK={lv_dlc_rotweak} SKY130_FD_PR__SPECIAL_NFET_LATCH__CDSC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__CDSCB_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__CDSCD_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__CIT_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__DLC_ROTWEAK={lv_dlc_rotweak} 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__DVT0_DIFF=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__DVT1_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__K2_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__K3_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__KT1_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__KT2_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__LINT_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__NFACTOR_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__TOX_SLOPE=0.005989 SKY130_FD_PR__SPECIAL_NFET_LATCH__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__VOFF_SLOPE=0.0 SKY130_FD_PR__SPECIAL_NFET_LATCH__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH__VTH0_SLOPE=0.005289 SKY130_FD_PR__SPECIAL_NFET_LATCH__WINT_SLOPE=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_LATCH_LOWLEAKAGE__DLC_ROTWEAK={lv_dlc_rotweak} SKY130_FD_PR__NFET_01V8__A0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_41=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_50=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_51=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_52=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_53=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_54=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_55=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_56=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_57=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_58=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_59=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_60=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_62=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8__A0_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_41=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_50=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_51=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_52=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_53=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_54=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_55=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_56=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_57=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_58=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_59=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_60=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_62=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__AGS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8__DLC_ROTWEAK={lv_dlc_rotweak} SKY130_FD_PR__NFET_01V8__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_40=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_42=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_44=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_46=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_48=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_49=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_50=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_62=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8__ETA0_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_38=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_41=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_50=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_51=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_56=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_57=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_58=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_59=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_60=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_61=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_62=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_40=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_42=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_44=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_46=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_48=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_49=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_50=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_52=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_53=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_54=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_55=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_59=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_60=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_62=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8__LINT_SLOPE=0.0 SKY130_FD_PR__NFET_01V8__NFACTOR_SLOPE=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_38=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_41=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_50=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_61=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_62=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8__PCLM_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_40=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_42=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_44=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_46=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_48=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_49=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_50=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_51=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_52=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_53=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_54=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_55=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_56=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_57=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_58=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_59=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_60=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_62=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_38=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_41=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_50=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_51=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_52=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_53=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_54=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_55=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_56=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_57=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_58=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_59=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_60=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_61=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_62=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8__PDITSD_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_40=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_42=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_43=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_44=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_45=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_46=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_47=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_48=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_49=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_50=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_51=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_52=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_53=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_54=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_55=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_56=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_57=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_58=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_59=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_60=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_61=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_62=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_01V8__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_01V8__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__RF_NFET_01V8__B_TOXE_SLOPE=0.003443 SKY130_FD_PR__RF_NFET_01V8__B_VOFF_SLOPE=0.007 
+ SKY130_FD_PR__RF_NFET_01V8__B_VTH0_SLOPE=0.005556 SKY130_FD_PR__RF_NFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8__BASE__DLC_ROTWEAK=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8__LINT1_SLOPE=0.0 
+ SKY130_FD_PR__RF_NFET_01V8__LINT_SLOPE=5.767e-9 SKY130_FD_PR__RF_NFET_01V8__TOXE1_SLOPE=0.006989 
+ SKY130_FD_PR__RF_NFET_01V8__TOXE2_SLOPE=0.005989 SKY130_FD_PR__RF_NFET_01V8__TOXE3_SLOPE=0.01089 
+ SKY130_FD_PR__RF_NFET_01V8__TOXE4_SLOPE=0.01289 SKY130_FD_PR__RF_NFET_01V8__TOXE_SLOPE=0.008989 
+ SKY130_FD_PR__NFET_01V8__RSHN_MULT=1.0 SKY130_FD_PR__NFET_01V8__TOXE_SLOPE=0.003443 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_11=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_12=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_13=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_14=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_15=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_16=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_17=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_18=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_19=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_20=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_21=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_22=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_23=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_24=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_25=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_26=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_27=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_28=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_29=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_30=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_31=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_32=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_33=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_34=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_35=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_36=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_37=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_38=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_39=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_40=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_41=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_42=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_50=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_51=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_52=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_53=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_54=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_55=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_56=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_57=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_58=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_59=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_60=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_61=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_62=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_15=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_16=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_17=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_18=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_23=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_24=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_25=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_26=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_31=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_32=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_33=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_34=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_40=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_41=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_47=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_48=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_49=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_50=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_51=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_52=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_53=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_54=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_55=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_56=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_57=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_58=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_59=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_60=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_61=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_62=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_01V8__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_01V8__VOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_01V8__VOFF_SLOPE=0.007 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_11=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_12=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_13=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_14=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_19=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_20=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_21=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_22=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_27=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_28=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_29=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_3=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_30=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_35=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_36=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_37=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_38=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_39=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_43=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_44=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_45=0.0 SKY130_FD_PR__NFET_01V8__VSAT_DIFF_46=0.0 
+ SKY130_FD_PR__NFET_01V8__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_01V8__VTH0_SLOPE=0.003356 
+ SKY130_FD_PR__NFET_01V8__VTH0_SLOPE1=0.007356 SKY130_FD_PR__NFET_01V8__WINT_SLOPE=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__AGS_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__B0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__B1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__B1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__DLC_ROTWEAK={lv_dlc_rotweak} SKY130_FD_PR__ESD_NFET_01V8__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__KETA_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__KETA_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PCLM_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PCLM_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITS_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITSD_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__PDITSD_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_01V8__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__RSHN_MULT=1.0 SKY130_FD_PR__ESD_NFET_01V8__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__TVOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_01V8__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__VOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_01V8__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_01V8__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__KU0_DIFF=-3.0e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__KVSAT_DIFF=0.3 SKY130_FD_PR__NFET_03V3_NVT__KVTH0_DIFF=-2.0e-9 
+ SKY130_FD_PR__NFET_03V3_NVT__LINT_SLOPE=0.0 SKY130_FD_PR__NFET_03V3_NVT__LKU0_DIFF=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__LKVTH0_DIFF=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_SLOPE=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RSHN_MULT=1.0 SKY130_FD_PR__NFET_03V3_NVT__TOXE_SLOPE=0.0045 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_SLOPE=0.0065 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_SLOPE=0.006 SKY130_FD_PR__NFET_03V3_NVT__WINT_SLOPE=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__WKU0_DIFF=5.0e-7 SKY130_FD_PR__NFET_03V3_NVT__WKVTH0_DIFF=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__WLOD_DIFF=0.0 SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KU0_DIFF=-9.9e-8 SKY130_FD_PR__NFET_G5V0D16V0__KVSAT_DIFF=0.3 
+ SKY130_FD_PR__NFET_G5V0D16V0__KVTH0_DIFF=1.7057e-8 SKY130_FD_PR__NFET_G5V0D16V0__LKU0_DIFF=9.6975e-7 
+ SKY130_FD_PR__NFET_G5V0D16V0__LKVTH0_DIFF=2.2691e-7 SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__WKU0_DIFF=2.0e-7 SKY130_FD_PR__NFET_G5V0D16V0__WKVTH0_DIFF=2.3093e-6 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__A0_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGIDL_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_66=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_67=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_HVT__AGS_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_55=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_56=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_HVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_55=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__B1_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_66=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_67=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_HVT__BGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_52=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_53=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_54=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_55=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_56=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_57=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_58=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_59=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_60=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_61=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_62=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_63=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_64=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_66=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_67=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_HVT__CGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__DLC_ROTWEAK={lvhvt_dlc_rotweak} SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_64=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_HVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KETA_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_66=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_HVT__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__LINT_SLOPE=0.0 SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_SLOPE=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_SLOPE1=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_64=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_66=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_67=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PCLM_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_64=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_66=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_67=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITS_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_64=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_66=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_67=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__PDITSD_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_64=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_66=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_67=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__RDSW_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__RSHP_MULT=1.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TOXE_SLOPE=0.005 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_52=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_53=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_54=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_55=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_59=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_60=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_61=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_62=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_63=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_64=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_65=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_66=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_67=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_HVT__UA_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__UA_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__UA_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__UA_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__UB_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__UB_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__UB_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__UB_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__VOFF_DIFF_56=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VOFF_DIFF_57=0.0 SKY130_FD_PR__PFET_01V8_HVT__VOFF_DIFF_58=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VOFF_DIFF_65=0.0 SKY130_FD_PR__PFET_01V8_HVT__VOFF_SLOPE=0.01 
+ SKY130_FD_PR__PFET_01V8_HVT__VOFF_SLOPE1=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8_HVT__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_HVT__VTH0_SLOPE=0.0055 SKY130_FD_PR__PFET_01V8_HVT__WINT_SLOPE=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_44=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__A0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGIDL_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_22=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_8=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_22=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_44=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_G5V0D10V5__BGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__ETA0_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_22=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_44=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_8=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KETA_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__KT1_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__KU0_DIFF=7.0e-8 
+ SKY130_FD_PR__PFET_G5V0D10V5__KVSAT_DIFF=0.4 SKY130_FD_PR__PFET_G5V0D10V5__KVTH0_DIFF=3.5e-8 
+ SKY130_FD_PR__PFET_G5V0D10V5__LINT_SLOPE=0.0 SKY130_FD_PR__PFET_G5V0D10V5__LKU0_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__LKVTH0_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D10V5__NFACTOR_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__NFACTOR_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__NFACTOR_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__NFACTOR_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__NFACTOR_SLOPE=0.02 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PCLM_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_22=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_44=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_8=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_27=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_29=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_30=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_32=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_34=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_38=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__PDITSD_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_22=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_44=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_8=0.0 SKY130_FD_PR__PFET_G5V0D10V5__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__RSHP_MULT=1.0 SKY130_FD_PR__PFET_G5V0D10V5__TOXE_SLOPE=0.012 
+ SKY130_FD_PR__PFET_G5V0D10V5__TOXE_SLOPE1=0.02 SKY130_FD_PR__PFET_G5V0D10V5__TOXE_SLOPE2=0.023 
+ SKY130_FD_PR__PFET_G5V0D10V5__TOXE_SLOPE3=0.014 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_11=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_13=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_15=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_20=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_22=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_40=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_42=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_44=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_46=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_48=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_8=0.0 SKY130_FD_PR__PFET_G5V0D10V5__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_10=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_12=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_16=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_18=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_21=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_24=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_26=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_28=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_33=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_36=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_41=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_47=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_5=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VOFF_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VOFF_SLOPE=0.009 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_14=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_17=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_19=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_23=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_25=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_3=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_31=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_35=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_37=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_39=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_43=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_45=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_7=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__VSAT_DIFF_9=0.0 SKY130_FD_PR__PFET_G5V0D10V5__VTH0_SLOPE=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__WINT_SLOPE=0.0 SKY130_FD_PR__PFET_G5V0D10V5__WKU0_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D10V5__WKVTH0_DIFF=6.5e-7 SKY130_FD_PR__PFET_G5V0D10V5__WLOD_DIFF=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__DLC_ROTWEAK={hv_dlc_rotweak} SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RSHP_MULT=1.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__A0_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__AGS_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B0_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__BGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__CGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__DLC_ROTWEAK={lvt_dlc_rotweak} SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__ETA0_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__KETA_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KU0_DIFF=5.9e-8 SKY130_FD_PR__PFET_01V8_LVT__KVSAT_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__KVTH0_DIFF=1.76e-8 SKY130_FD_PR__PFET_01V8_LVT__LINT_SLOPE=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__LKU0_DIFF=0.0 SKY130_FD_PR__PFET_01V8_LVT__LKVTH0_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_SLOPE=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PCLM_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITS_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__PDITSD_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RDSW_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__RF_BASE_DLC_ROTWEAK=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__RSHP_MULT=1.0 SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE=0.003689 
+ SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE1=0.01489 SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE2=0.01689 
+ SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE3=0.02389 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UA_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__UB_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VOFF_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8_LVT__VOFF_SLOPE=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8_LVT__VSAT_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE=0.01389 SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE1=0.009789 
+ SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE2=0.01089 SKY130_FD_PR__PFET_01V8_LVT__WINT_SLOPE=0.0 
+ SKY130_FD_PR__PFET_01V8_LVT__WKU0_DIFF=0.0 SKY130_FD_PR__PFET_01V8_LVT__WKVTH0_DIFF=7.3e-7 
+ SKY130_FD_PR__PFET_01V8_LVT__WLOD_DIFF=0.0 SKY130_FD_PR__PFET_01V8_MVT__A0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__A0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__AGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__AGS_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__B0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__B1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__BGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__CGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__KT1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8_MVT__NFACTOR_SLOPE=0.1 
+ SKY130_FD_PR__PFET_01V8_MVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__PDITSD_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RD_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_MVT__AW_RS_MULT=1.0 
+ SKY130_FD_PR__PFET_01V8_MVT__RSHP_MULT=1.0 SKY130_FD_PR__PFET_01V8_MVT__TOXE_SLOPE=0.025 
+ SKY130_FD_PR__PFET_01V8_MVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__UA_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__UA_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__UB_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__UB_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__VOFF_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8_MVT__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8_MVT__VOFF_SLOPE=0.0 SKY130_FD_PR__PFET_01V8_MVT__VTH0_SLOPE=0.05 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__CDSC_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__CDSCB_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__CDSCD_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__CIT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__DLC_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__DLC_ROTWEAK={lv_dlc_rotweak} 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__DVT0_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__DWC_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__K2_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__K3_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__KT1_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__KT1L_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__KT2_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__LINT_DIFF=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__LINT_SLOPE=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__NFACTOR_SLOPE=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__TOX_MULT=1.0 SKY130_FD_PR__SPECIAL_PFET_PASS__TOX_SLOPE=0.005567 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__VOFF_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__VOFF_SLOPE=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__VSAT_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__VTH0_SLOPE=0.005567 
+ SKY130_FD_PR__SPECIAL_PFET_PASS__WINT_DIFF=0.0 SKY130_FD_PR__SPECIAL_PFET_PASS__WINT_SLOPE=0.0 
+ SKY130_FD_PR__SPECIAL_PFET_PASS_LOWLEAKAGE__DLC_ROTWEAK={lv_dlc_rotweak} SKY130_FD_PR__PFET_01V8__A0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8__A0_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__A0_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__AGS_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__AGS_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8__B0_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__B0_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8__B1_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__B1_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__BGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__CGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__DLC_ROTWEAK={lv_dlc_rotweak} SKY130_FD_PR__PFET_01V8__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8__ETA0_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8__KETA_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_1=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_11=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_15=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_16=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_17=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_18=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_23=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_24=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_25=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_26=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_31=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_32=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_33=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_34=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_36=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_37=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_38=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_39=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_40=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_41=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_42=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_43=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_45=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_46=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_47=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_48=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_49=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_50=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_51=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_7=0.0 SKY130_FD_PR__PFET_01V8__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__PFET_01V8__KT1_DIFF_9=0.0 SKY130_FD_PR__PFET_01V8__KU0_DIFF=4.5e-8 
+ SKY130_FD_PR__PFET_01V8__KVSAT_DIFF=0.5 SKY130_FD_PR__PFET_01V8__KVTH0_DIFF=3.29e-8 
+ SKY130_FD_PR__PFET_01V8__LINT_SLOPE=0.0 SKY130_FD_PR__PFET_01V8__LKU0_DIFF=0.0 
+ SKY130_FD_PR__PFET_01V8__LKVTH0_DIFF=0.0 SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE=0.1 
+ SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE1=0.1 SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE2=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__PCLM_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITS_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__RDSW_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RD_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8__AW_RS_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__B_NFACTOR_SLOPE1=0.1 SKY130_FD_PR__RF_PFET_01V8__B_TOXE_SLOPE=0.006443 
+ SKY130_FD_PR__RF_PFET_01V8__B_TOXE_SLOPE1=0.004443 SKY130_FD_PR__RF_PFET_01V8__B_VOFF_SLOPE=0.014 
+ SKY130_FD_PR__RF_PFET_01V8__B_VOFF_SLOPE1=0.009 SKY130_FD_PR__RF_PFET_01V8__B_VTH0_SLOPE1=0.007356 
+ SKY130_FD_PR__RF_PFET_01V8__B_VTH0_SLOPE2=0.009356 SKY130_FD_PR__RF_PFET_01V8__B_VTH0_SLOPE3=0.008356 
+ SKY130_FD_PR__RF_PFET_01V8_B__DWC_DIFF=0.0 SKY130_FD_PR__RF_PFET_01V8__BASE__DLC_ROTWEAK=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8__NFACTOR1_SLOPE=0.0 SKY130_FD_PR__RF_PFET_01V8__NFACTOR_SLOPE=0.429 
+ SKY130_FD_PR__RF_PFET_01V8__TOXE1_SLOPE=0.01067 SKY130_FD_PR__RF_PFET_01V8__TOXE2_SLOPE=0.01167 
+ SKY130_FD_PR__RF_PFET_01V8__TOXE3_SLOPE=0.01367 SKY130_FD_PR__RF_PFET_01V8__TOXE4_SLOPE=0.01467 
+ SKY130_FD_PR__RF_PFET_01V8__TOXE5_SLOPE=0.01567 SKY130_FD_PR__RF_PFET_01V8__TOXE_SLOPE=0.01267 
+ SKY130_FD_PR__PFET_01V8__RSHP_MULT=1.0 SKY130_FD_PR__PFET_01V8__TOXE_SLOPE=0.004443 
+ SKY130_FD_PR__PFET_01V8__TOXE_SLOPE1=0.006443 SKY130_FD_PR__PFET_01V8__TOXE_SLOPE2=0.003443 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_0=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_10=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_11=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_12=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_13=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_14=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_15=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_16=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_17=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_18=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_19=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_2=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_20=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_21=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_22=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_23=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_24=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_25=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_26=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_27=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_28=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_29=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_30=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_31=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_32=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_33=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_34=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_35=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_36=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_39=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_4=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_40=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_41=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_42=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_43=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_44=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_45=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_47=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_48=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_49=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_50=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_51=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_6=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_8=0.0 SKY130_FD_PR__PFET_01V8__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__PFET_01V8__VOFF_SLOPE=0.0 SKY130_FD_PR__PFET_01V8__VOFF_SLOPE1=0.0 
+ SKY130_FD_PR__PFET_01V8__VOFF_SLOPE2=0.007 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_12=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_13=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_14=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_19=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_20=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_21=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_22=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_27=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_28=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_29=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_3=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_30=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_35=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_37=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_38=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_44=0.0 SKY130_FD_PR__PFET_01V8__VSAT_DIFF_46=0.0 
+ SKY130_FD_PR__PFET_01V8__VSAT_DIFF_5=0.0 SKY130_FD_PR__PFET_01V8__VTH0_SLOPE=0.005856 
+ SKY130_FD_PR__PFET_01V8__VTH0_SLOPE1=0.007356 SKY130_FD_PR__PFET_01V8__VTH0_SLOPE2=0.004356 
+ SKY130_FD_PR__PFET_01V8__WINT_SLOPE=0.0 SKY130_FD_PR__PFET_01V8__WKU0_DIFF=2.5e-7 
+ SKY130_FD_PR__PFET_01V8__WKVTH0_DIFF=2.0e-7 SKY130_FD_PR__PFET_01V8__WLOD_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__A0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__A0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AGS_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGBACC_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGBACC_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGBINV_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGBINV_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGC_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGC_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGSD_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__B0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__B0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__B1_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__B1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__BGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__BIGSD_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__BIGSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__CF_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D16V0__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__CGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__CJSWGS_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__DLC_ROTWEAK={hv_dlc_rotweak} SKY130_FD_PR__PFET_G5V0D16V0__DSUB_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__DSUB_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__ETA0_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__JTSSWS_DIFF_0=-4.02e-12 
+ SKY130_FD_PR__PFET_G5V0D16V0__JTSSWS_DIFF_1=-4.02e-12 SKY130_FD_PR__PFET_G5V0D16V0__K2_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__K2_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__KT1_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__KU0_DIFF=2.218e-7 
+ SKY130_FD_PR__PFET_G5V0D16V0__KVSAT_DIFF=0.4 SKY130_FD_PR__PFET_G5V0D16V0__KVTH0_DIFF=5.2302e-9 
+ SKY130_FD_PR__PFET_G5V0D16V0__LKU0_DIFF=8.7129e-7 SKY130_FD_PR__PFET_G5V0D16V0__LKVTH0_DIFF=-4.8631e-7 
+ SKY130_FD_PR__PFET_G5V0D16V0__LPE0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__LPE0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__NIGBACC_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__NIGBACC_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__NIGBINV_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__NIGBINV_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PCLM_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PDITS_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PDITSD_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__RDSW_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__RDW_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__RDW_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__RSHP_MULT=1.0 SKY130_FD_PR__PFET_G5V0D16V0__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__TVOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__UA_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__UA_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__UB_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__UB_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VSAT_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__WKU0_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__WKVTH0_DIFF=5.398e-7 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__AJUNCTION_MULT=1.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__DLC_DIFF=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__DWC_DIFF=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__K2_DIFF_0=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__K2_DIFF_1=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__K2_DIFF_2=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__KT1_DIFF_0=-0.44275 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__KT1_DIFF_1=-0.3267 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__KT1_DIFF_2=-0.67944 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__LINT_DIFF=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__NFACTOR_DIFF_0=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__NFACTOR_DIFF_2=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__OVERLAP_MULT=1.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__PJUNCTION_MULT=1.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__RDSW_DIFF_0=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__RDSW_DIFF_1=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__RDSW_DIFF_2=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__TOX_MULT=1.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__TOX_SLOPE=0.002 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__TOX_SLOPE1=0.002 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__U0_DIFF_0=-0.0069221 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__U0_DIFF_1=-0.0041919 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__U0_DIFF_2=-0.0081788 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VOFF_DIFF_0=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VOFF_DIFF_1=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VOFF_DIFF_2=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VSAT_DIFF_0=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VSAT_DIFF_1=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VSAT_DIFF_2=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_DIFF_0=0.91203 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_DIFF_1=1.3659 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_DIFF_2=0.27494 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_SLOPE=0.0255 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_SLOPE1=0.028 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__WINT_DIFF=0.0 
+ SONOS_EEOL_DLC_ROTWEAK={hv_dlc_rotweak} SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__AJUNCTION_MULT=1.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__DLC_DIFF=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__DLC_ROTWEAK={hv_dlc_rotweak} 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__DWC_DIFF=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__K2_DIFF_0=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__K2_DIFF_1=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__K2_DIFF_2=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__KT1_DIFF_0=-0.36466 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__KT1_DIFF_1=-0.029107 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__KT1_DIFF_2=-0.65907 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__LINT_DIFF=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__NFACTOR_DIFF_0=-0.23845 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__NFACTOR_DIFF_1=1.3597 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__NFACTOR_DIFF_2=1.0202 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__OVERLAP_MULT=1.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__PJUNCTION_MULT=1.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__RDSW_DIFF_0=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__RDSW_DIFF_1=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__RDSW_DIFF_2=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__TOX_MULT=1.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__TOX_SLOPE=0.005 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__U0_DIFF_0=-0.004 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__U0_DIFF_1=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__U0_DIFF_2=0.0013468 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VOFF_DIFF_0=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VOFF_DIFF_1=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VOFF_DIFF_2=-0.20912 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VSAT_DIFF_0=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VSAT_DIFF_1=0.0 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VSAT_DIFF_2=0.0 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VTH0_DIFF_0=-1.0278 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VTH0_DIFF_1=-0.85561 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VTH0_DIFF_2=-0.15565 
+ SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__VTH0_SLOPE=0.026 SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_ORIGINAL__WINT_DIFF=0.0 
+ SONOS_PEOL_DLC_ROTWEAK={hv_dlc_rotweak} SKY130_FD_PR__NFET_20V0_NVT__REVERSE_TMAX='20.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT__REVERSE_VDS='-0.01' SKY130_FD_PR__NFET_20V0_NVT__TMAX_VBD_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT__TMAX_VBD_2='25.001n' SKY130_FD_PR__NFET_20V0_NVT__TMAX_VBS_1='20.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT__TMAX_VDS_1='100.001n' SKY130_FD_PR__NFET_20V0_NVT__TMAX_VDS_2='25.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT__TMAX_VGB_1='100.001n' SKY130_FD_PR__NFET_20V0_NVT__TMAX_VGB_2='20.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT__TMAX_VGD_1='sky130_fd_pr__nfet_20v0_nvt__tmax_vds_1' 
+ SKY130_FD_PR__NFET_20V0_NVT__TMAX_VGD_2='sky130_fd_pr__nfet_20v0_nvt__tmax_vds_2' 
+ SKY130_FD_PR__NFET_20V0_NVT__TMAX_VGS_1='100.001n' SKY130_FD_PR__NFET_20V0_NVT__TMAX_VGS_2='20.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBD_MAX='sky130_fd_pr__nfet_20v0_nvt__vbs_max' SKY130_FD_PR__NFET_20V0_NVT__VBD_MAX_1='sky130_fd_pr__nfet_20v0_nvt__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBD_MAX_2='sky130_fd_pr__nfet_20v0_nvt__vbs_max' SKY130_FD_PR__NFET_20V0_NVT__VBD_MIN='sky130_fd_pr__nfet_20v0_nvt__vbs_min - sky130_fd_pr__nfet_20v0_nvt__vds_max' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBD_MIN_1='sky130_fd_pr__nfet_20v0_nvt__vbs_min - sky130_fd_pr__nfet_20v0_nvt__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBD_MIN_2='sky130_fd_pr__nfet_20v0_nvt__vbs_min - sky130_fd_pr__nfet_20v0_nvt__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBD_REVERSEMAX='0.501' SKY130_FD_PR__NFET_20V0_NVT__VBD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBS_MAX='0.001' SKY130_FD_PR__NFET_20V0_NVT__VBS_MAX_1='0.001' 
+ SKY130_FD_PR__NFET_20V0_NVT__VBS_MIN='-2.501' SKY130_FD_PR__NFET_20V0_NVT__VBS_MIN_1='-2.501' 
+ SKY130_FD_PR__NFET_20V0_NVT__VDS_MAX='36' SKY130_FD_PR__NFET_20V0_NVT__VDS_MAX_1='24.501' 
+ SKY130_FD_PR__NFET_20V0_NVT__VDS_MAX_2='30.001' SKY130_FD_PR__NFET_20V0_NVT__VDS_MIN='-0.001' 
+ SKY130_FD_PR__NFET_20V0_NVT__VDS_MIN_1='-0.001' SKY130_FD_PR__NFET_20V0_NVT__VDS_MIN_2='-0.001' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGB_MAX='sky130_fd_pr__nfet_20v0_nvt__vgs_max - sky130_fd_pr__nfet_20v0_nvt__vbs_min' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGB_MAX_1='sky130_fd_pr__nfet_20v0_nvt__vgs_max_1 - sky130_fd_pr__nfet_20v0_nvt__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGB_MAX_2='sky130_fd_pr__nfet_20v0_nvt__vgs_max_2 - sky130_fd_pr__nfet_20v0_nvt__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGB_MIN='-1*sky130_fd_pr__nfet_20v0_nvt__vgs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGB_MIN_1='0 - 2.5' SKY130_FD_PR__NFET_20V0_NVT__VGB_MIN_2='0 - 2.5' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_MAX='sky130_fd_pr__nfet_20v0_nvt__vgs_max' SKY130_FD_PR__NFET_20V0_NVT__VGD_MAX_1='sky130_fd_pr__nfet_20v0_nvt__vgs_max_1' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_MAX_2='sky130_fd_pr__nfet_20v0_nvt__vgs_max_2' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_MIN='-1*sky130_fd_pr__nfet_20v0_nvt__vds_max' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_MIN_1='-1*sky130_fd_pr__nfet_20v0_nvt__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_MIN_2='-1*sky130_fd_pr__nfet_20v0_nvt__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_NVT__VGD_REVERSEMAX_1='0.101' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGD_REVERSEMIN='-5.501' SKY130_FD_PR__NFET_20V0_NVT__VGD_REVERSEMIN_1='-0.101' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGS_MAX='6.501' SKY130_FD_PR__NFET_20V0_NVT__VGS_MAX_1='5.751' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGS_MAX_2='6.001' SKY130_FD_PR__NFET_20V0_NVT__VGS_MIN='-1*6.501' 
+ SKY130_FD_PR__NFET_20V0_NVT__VGS_MIN_1='-1*5.751' SKY130_FD_PR__NFET_20V0_NVT__VGS_MIN_2='-1*6.001' 
+ SKY130_FD_PR__NFET_20V0_NVT__VSD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_NVT__VSD_REVERSEMIN='-0.501' 
+ SKY130_FD_PR__NFET_20V0_NVT__VTX='0.020' SKY130_FD_PR__NFET_20V0_NVT_ISO__K2_DIFF=-0.11937 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__REVERSE_TMAX='20.001n' SKY130_FD_PR__NFET_20V0_NVT_ISO__REVERSE_VDS='-0.01' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VBD_1='100.001n' SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VBD_2='25.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VBS_1='20.001n' SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VDS_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VDS_2='25.001n' SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VGB_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VGB_2='20.001n' SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VGD_1='sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_1' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VGD_2='sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_2' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VGS_1='100.001n' SKY130_FD_PR__NFET_20V0_NVT_ISO__TMAX_VGS_2='20.001n' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_MAX='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_MAX_1='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_MAX_2='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_MIN='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min - sky130_fd_pr__nfet_20v0_nvt_iso__vds_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_MIN_1='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min - sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_MIN_2='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min - sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_REVERSEMAX='0.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VBD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBS_MAX='0.001' SKY130_FD_PR__NFET_20V0_NVT_ISO__VBS_MAX_1='0.001' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VBS_MIN='-2.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VBS_MIN_1='-2.501' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VDS_MAX='22.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VDS_MAX_1='22.001' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VDS_MAX_2='22.001' SKY130_FD_PR__NFET_20V0_NVT_ISO__VDS_MIN='-0.001' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VDS_MIN_1='-0.001' SKY130_FD_PR__NFET_20V0_NVT_ISO__VDS_MIN_2='-0.001' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGB_MAX='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max - sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGB_MAX_1='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1 - sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGB_MAX_2='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2 - sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGB_MIN='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGB_MIN_1='0 - 2.5' SKY130_FD_PR__NFET_20V0_NVT_ISO__VGB_MIN_2='0 - 2.5' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_MAX='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_MAX_1='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_MAX_2='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_MIN='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_MIN_1='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_MIN_2='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_REVERSEMAX_1='0.101' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_REVERSEMIN='-5.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VGD_REVERSEMIN_1='-0.101' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGS_MAX='6.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VGS_MAX_1='5.751' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGS_MAX_2='6.001' SKY130_FD_PR__NFET_20V0_NVT_ISO__VGS_MIN='-1*6.501' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VGS_MIN_1='-1*5.751' SKY130_FD_PR__NFET_20V0_NVT_ISO__VGS_MIN_2='-1*6.001' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VSD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_NVT_ISO__VSD_REVERSEMIN='-0.501' 
+ SKY130_FD_PR__NFET_20V0_NVT_ISO__VTX='0.02' SKY130_FD_PR__NFET_20V0__REVERSE_TMAX='20.001n' 
+ SKY130_FD_PR__NFET_20V0__REVERSE_VDS='-0.01' SKY130_FD_PR__NFET_20V0__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_20V0__TMAX_VBD_1='100.001n' SKY130_FD_PR__NFET_20V0__TMAX_VBD_2='25.001n' 
+ SKY130_FD_PR__NFET_20V0__TMAX_VBS_1='20.001n' SKY130_FD_PR__NFET_20V0__TMAX_VDS_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0__TMAX_VDS_2='25.001n' SKY130_FD_PR__NFET_20V0__TMAX_VGB_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0__TMAX_VGB_2='20.001n' SKY130_FD_PR__NFET_20V0__TMAX_VGD_1='sky130_fd_pr__nfet_20v0__tmax_vds_1' 
+ SKY130_FD_PR__NFET_20V0__TMAX_VGD_2='sky130_fd_pr__nfet_20v0__tmax_vds_2' SKY130_FD_PR__NFET_20V0__TMAX_VGS_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0__TMAX_VGS_2='20.001n' SKY130_FD_PR__NFET_20V0__VBD_MAX='sky130_fd_pr__nfet_20v0__vbs_max' 
+ SKY130_FD_PR__NFET_20V0__VBD_MAX_1='sky130_fd_pr__nfet_20v0__vbs_max' SKY130_FD_PR__NFET_20V0__VBD_MAX_2='sky130_fd_pr__nfet_20v0__vbs_max' 
+ SKY130_FD_PR__NFET_20V0__VBD_MIN='sky130_fd_pr__nfet_20v0__vbs_min - sky130_fd_pr__nfet_20v0__vds_max' 
+ SKY130_FD_PR__NFET_20V0__VBD_MIN_1='sky130_fd_pr__nfet_20v0__vbs_min - sky130_fd_pr__nfet_20v0__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0__VBD_MIN_2='sky130_fd_pr__nfet_20v0__vbs_min - sky130_fd_pr__nfet_20v0__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0__VBD_REVERSEMAX='0.501' SKY130_FD_PR__NFET_20V0__VBD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__NFET_20V0__VBS_MAX='0.001' SKY130_FD_PR__NFET_20V0__VBS_MAX_1='0.001' 
+ SKY130_FD_PR__NFET_20V0__VBS_MIN='-2.501' SKY130_FD_PR__NFET_20V0__VBS_MIN_1='-2.501' 
+ SKY130_FD_PR__NFET_20V0__VDS_MAX='36' SKY130_FD_PR__NFET_20V0__VDS_MAX_1='24.501' 
+ SKY130_FD_PR__NFET_20V0__VDS_MAX_2='30.001' SKY130_FD_PR__NFET_20V0__VDS_MIN='-0.001' 
+ SKY130_FD_PR__NFET_20V0__VDS_MIN_1='-0.001' SKY130_FD_PR__NFET_20V0__VDS_MIN_2='-0.001' 
+ SKY130_FD_PR__NFET_20V0__VGB_MAX='sky130_fd_pr__nfet_20v0__vgs_max - sky130_fd_pr__nfet_20v0__vbs_min' 
+ SKY130_FD_PR__NFET_20V0__VGB_MAX_1='sky130_fd_pr__nfet_20v0__vgs_max_1 - sky130_fd_pr__nfet_20v0__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0__VGB_MAX_2='sky130_fd_pr__nfet_20v0__vgs_max_2 - sky130_fd_pr__nfet_20v0__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0__VGB_MIN='-1*sky130_fd_pr__nfet_20v0__vgs_max' SKY130_FD_PR__NFET_20V0__VGB_MIN_1='0 - 2.5' 
+ SKY130_FD_PR__NFET_20V0__VGB_MIN_2='0 - 2.5' SKY130_FD_PR__NFET_20V0__VGD_MAX='sky130_fd_pr__nfet_20v0__vgs_max' 
+ SKY130_FD_PR__NFET_20V0__VGD_MAX_1='sky130_fd_pr__nfet_20v0__vgs_max_1' SKY130_FD_PR__NFET_20V0__VGD_MAX_2='sky130_fd_pr__nfet_20v0__vgs_max_2' 
+ SKY130_FD_PR__NFET_20V0__VGD_MIN='-1*sky130_fd_pr__nfet_20v0__vds_max' SKY130_FD_PR__NFET_20V0__VGD_MIN_1='-1*sky130_fd_pr__nfet_20v0__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0__VGD_MIN_2='-1*sky130_fd_pr__nfet_20v0__vds_max_2' SKY130_FD_PR__NFET_20V0__VGD_REVERSEMAX='5.501' 
+ SKY130_FD_PR__NFET_20V0__VGD_REVERSEMAX_1='0.101' SKY130_FD_PR__NFET_20V0__VGD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__NFET_20V0__VGD_REVERSEMIN_1='-0.101' SKY130_FD_PR__NFET_20V0__VGS_MAX='6.501' 
+ SKY130_FD_PR__NFET_20V0__VGS_MAX_1='5.751' SKY130_FD_PR__NFET_20V0__VGS_MAX_2='6.001' 
+ SKY130_FD_PR__NFET_20V0__VGS_MIN='-1*6.501' SKY130_FD_PR__NFET_20V0__VGS_MIN_1='-1*5.751' 
+ SKY130_FD_PR__NFET_20V0__VGS_MIN_2='-1*6.001' SKY130_FD_PR__NFET_20V0__VSD_REVERSEMAX='5.501' 
+ SKY130_FD_PR__NFET_20V0__VSD_REVERSEMIN='-0.501' SKY130_FD_PR__NFET_20V0__VTX='0.623' 
+ SKY130_FD_PR__NFET_20V0_ISO__REVERSE_TMAX='20.001n' SKY130_FD_PR__NFET_20V0_ISO__REVERSE_VDS='-0.01' 
+ SKY130_FD_PR__NFET_20V0_ISO__TMAX_VBD_1='100.001n' SKY130_FD_PR__NFET_20V0_ISO__TMAX_VBD_2='25.001n' 
+ SKY130_FD_PR__NFET_20V0_ISO__TMAX_VBS_1='20.001n' SKY130_FD_PR__NFET_20V0_ISO__TMAX_VDS_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_ISO__TMAX_VDS_2='25.001n' SKY130_FD_PR__NFET_20V0_ISO__TMAX_VGB_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_ISO__TMAX_VGB_2='20.001n' SKY130_FD_PR__NFET_20V0_ISO__TMAX_VGD_1='sky130_fd_pr__nfet_20v0_iso__tmax_vds_1' 
+ SKY130_FD_PR__NFET_20V0_ISO__TMAX_VGD_2='sky130_fd_pr__nfet_20v0_iso__tmax_vds_2' 
+ SKY130_FD_PR__NFET_20V0_ISO__TMAX_VGS_1='100.001n' SKY130_FD_PR__NFET_20V0_ISO__TMAX_VGS_2='20.001n' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBD_MAX='sky130_fd_pr__nfet_20v0_iso__vbs_max' SKY130_FD_PR__NFET_20V0_ISO__VBD_MAX_1='sky130_fd_pr__nfet_20v0_iso__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBD_MAX_2='sky130_fd_pr__nfet_20v0_iso__vbs_max' SKY130_FD_PR__NFET_20V0_ISO__VBD_MIN='sky130_fd_pr__nfet_20v0_iso__vbs_min - sky130_fd_pr__nfet_20v0_iso__vds_max' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBD_MIN_1='sky130_fd_pr__nfet_20v0_iso__vbs_min - sky130_fd_pr__nfet_20v0_iso__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBD_MIN_2='sky130_fd_pr__nfet_20v0_iso__vbs_min - sky130_fd_pr__nfet_20v0_iso__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBD_REVERSEMAX='0.501' SKY130_FD_PR__NFET_20V0_ISO__VBD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBS_MAX='0.001' SKY130_FD_PR__NFET_20V0_ISO__VBS_MAX_1='0.001' 
+ SKY130_FD_PR__NFET_20V0_ISO__VBS_MIN='-2.501' SKY130_FD_PR__NFET_20V0_ISO__VBS_MIN_1='-2.501' 
+ SKY130_FD_PR__NFET_20V0_ISO__VDS_MAX='22.501' SKY130_FD_PR__NFET_20V0_ISO__VDS_MAX_1='22.001' 
+ SKY130_FD_PR__NFET_20V0_ISO__VDS_MAX_2='22.001' SKY130_FD_PR__NFET_20V0_ISO__VDS_MIN='-0.001' 
+ SKY130_FD_PR__NFET_20V0_ISO__VDS_MIN_1='-0.001' SKY130_FD_PR__NFET_20V0_ISO__VDS_MIN_2='-0.001' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGB_MAX='sky130_fd_pr__nfet_20v0_iso__vgs_max - sky130_fd_pr__nfet_20v0_iso__vbs_min' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGB_MAX_1='sky130_fd_pr__nfet_20v0_iso__vgs_max_1 - sky130_fd_pr__nfet_20v0_iso__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGB_MAX_2='sky130_fd_pr__nfet_20v0_iso__vgs_max_2 - sky130_fd_pr__nfet_20v0_iso__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGB_MIN='-1*sky130_fd_pr__nfet_20v0_iso__vgs_max' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGB_MIN_1='0 - 2.5' SKY130_FD_PR__NFET_20V0_ISO__VGB_MIN_2='0 - 2.5' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_MAX='sky130_fd_pr__nfet_20v0_iso__vgs_max' SKY130_FD_PR__NFET_20V0_ISO__VGD_MAX_1='sky130_fd_pr__nfet_20v0_iso__vgs_max_1' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_MAX_2='sky130_fd_pr__nfet_20v0_iso__vgs_max_2' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_MIN='-1*sky130_fd_pr__nfet_20v0_iso__vds_max' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_MIN_1='-1*sky130_fd_pr__nfet_20v0_iso__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_MIN_2='-1*sky130_fd_pr__nfet_20v0_iso__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_ISO__VGD_REVERSEMAX_1='0.101' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGD_REVERSEMIN='-5.501' SKY130_FD_PR__NFET_20V0_ISO__VGD_REVERSEMIN_1='-0.101' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGS_MAX='6.501' SKY130_FD_PR__NFET_20V0_ISO__VGS_MAX_1='5.751' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGS_MAX_2='6.001' SKY130_FD_PR__NFET_20V0_ISO__VGS_MIN='-1*6.501' 
+ SKY130_FD_PR__NFET_20V0_ISO__VGS_MIN_1='-1*5.751' SKY130_FD_PR__NFET_20V0_ISO__VGS_MIN_2='-1*6.001' 
+ SKY130_FD_PR__NFET_20V0_ISO__VSD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_ISO__VSD_REVERSEMIN='-0.501' 
+ SKY130_FD_PR__NFET_20V0_ISO__VTX='0.617' SKY130_FD_PR__NFET_20V0_ZVT__HVVSAT_MULT=1.0 
+ SKY130_FD_PR__NFET_20V0_ZVT__K2_DIFF=0.0 SKY130_FD_PR__NFET_20V0_ZVT__LINT_DIFF=0.0 
+ SKY130_FD_PR__NFET_20V0_ZVT__REVERSE_TMAX='20.001n' SKY130_FD_PR__NFET_20V0_ZVT__REVERSE_VDS='-0.01' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VBD_1='100.001n' SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VBD_2='25.001n' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VBS_1='20.001n' SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VDS_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VDS_2='25.001n' SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGB_1='100.001n' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGB_2='20.001n' SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGD_1='sky130_fd_pr__nfet_20v0_zvt__tmax_vds_1' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGD_2='sky130_fd_pr__nfet_20v0_zvt__tmax_vds_2' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGS_1='100.001n' SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGS_2='20.001n' 
+ SKY130_FD_PR__NFET_20V0_ZVT__TMAX_VGS_MODEL01='0.001n' SKY130_FD_PR__NFET_20V0_ZVT__VBD_MAX='sky130_fd_pr__nfet_20v0_zvt__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBD_MAX_1='sky130_fd_pr__nfet_20v0_zvt__vbs_max' SKY130_FD_PR__NFET_20V0_ZVT__VBD_MAX_2='sky130_fd_pr__nfet_20v0_zvt__vbs_max' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBD_MIN='sky130_fd_pr__nfet_20v0_zvt__vbs_min - sky130_fd_pr__nfet_20v0_zvt__vds_max' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBD_MIN_1='sky130_fd_pr__nfet_20v0_zvt__vbs_min - sky130_fd_pr__nfet_20v0_zvt__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBD_MIN_2='sky130_fd_pr__nfet_20v0_zvt__vbs_min - sky130_fd_pr__nfet_20v0_zvt__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBD_REVERSEMAX='0.501' SKY130_FD_PR__NFET_20V0_ZVT__VBD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBS_MAX='0.001' SKY130_FD_PR__NFET_20V0_ZVT__VBS_MAX_1='0.001' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VBS_MIN='-2.501' SKY130_FD_PR__NFET_20V0_ZVT__VBS_MIN_1='-2.501' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VDS_MAX='30.001' SKY130_FD_PR__NFET_20V0_ZVT__VDS_MAX_1='24.501' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VDS_MAX_2='28.001' SKY130_FD_PR__NFET_20V0_ZVT__VDS_MAX_MODEL01='1*3.0' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VDS_MIN='-0.001' SKY130_FD_PR__NFET_20V0_ZVT__VDS_MIN_1='-0.001' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VDS_MIN_2='-0.001' SKY130_FD_PR__NFET_20V0_ZVT__VDS_MIN_MODEL01='-1*3.0' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGB_MAX='sky130_fd_pr__nfet_20v0_zvt__vgs_max - sky130_fd_pr__nfet_20v0_zvt__vbs_min' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGB_MAX_1='sky130_fd_pr__nfet_20v0_zvt__vgs_max_1 - sky130_fd_pr__nfet_20v0_zvt__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGB_MAX_2='sky130_fd_pr__nfet_20v0_zvt__vgs_max_2 - sky130_fd_pr__nfet_20v0_zvt__vbs_min_1' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGB_MIN='-1*sky130_fd_pr__nfet_20v0_zvt__vgs_max' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGB_MIN_1='0 - 2.5' SKY130_FD_PR__NFET_20V0_ZVT__VGB_MIN_2='0 - 2.5' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_MAX='sky130_fd_pr__nfet_20v0_zvt__vgs_max' SKY130_FD_PR__NFET_20V0_ZVT__VGD_MAX_1='sky130_fd_pr__nfet_20v0_zvt__vgs_max_1' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_MAX_2='sky130_fd_pr__nfet_20v0_zvt__vgs_max_2' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_MIN='-1*sky130_fd_pr__nfet_20v0_zvt__vds_max' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_MIN_1='-1*sky130_fd_pr__nfet_20v0_zvt__vds_max_1' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_MIN_2='-1*sky130_fd_pr__nfet_20v0_zvt__vds_max_2' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_REVERSEMAX='5.501' SKY130_FD_PR__NFET_20V0_ZVT__VGD_REVERSEMAX_1='0.101' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGD_REVERSEMIN='-5.501' SKY130_FD_PR__NFET_20V0_ZVT__VGD_REVERSEMIN_1='-0.101' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGS_MAX='6.501' SKY130_FD_PR__NFET_20V0_ZVT__VGS_MAX_1='5.751' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGS_MAX_2='6.001' SKY130_FD_PR__NFET_20V0_ZVT__VGS_MAX_MODEL01='1*3.0' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGS_MIN='-1*6.501' SKY130_FD_PR__NFET_20V0_ZVT__VGS_MIN_1='-1*5.751' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGS_MIN_2='-1*6.001' SKY130_FD_PR__NFET_20V0_ZVT__VGS_MIN_MODEL01='-1*3.0' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VSAT_DIFF=0.0 SKY130_FD_PR__NFET_20V0_ZVT__VSD_REVERSEMAX='5.501' 
+ SKY130_FD_PR__NFET_20V0_ZVT__VSD_REVERSEMIN='-0.501' SKY130_FD_PR__NFET_20V0_ZVT__VTX='-0.223' 
+ SKY130_FD_PR__PFET_20V0__AGIDL_DIFF=0.0 SKY130_FD_PR__PFET_20V0__K2_DIFF=0.0 SKY130_FD_PR__PFET_20V0__REVERSE_TMAX='20.001n' 
+ SKY130_FD_PR__PFET_20V0__REVERSE_VDS='0.01' SKY130_FD_PR__PFET_20V0__RSHN_MULT=1.0 
+ SKY130_FD_PR__PFET_20V0__TMAX_VBD_1='100.001n' SKY130_FD_PR__PFET_20V0__TMAX_VBD_2='25.001n' 
+ SKY130_FD_PR__PFET_20V0__TMAX_VBS_1='20.001n' SKY130_FD_PR__PFET_20V0__TMAX_VDS_1='100.001n' 
+ SKY130_FD_PR__PFET_20V0__TMAX_VDS_2='25.001n' SKY130_FD_PR__PFET_20V0__TMAX_VGB_1='100.001n' 
+ SKY130_FD_PR__PFET_20V0__TMAX_VGB_2='20.001n' SKY130_FD_PR__PFET_20V0__TMAX_VGD_1='sky130_fd_pr__pfet_20v0__tmax_vds_1' 
+ SKY130_FD_PR__PFET_20V0__TMAX_VGD_2='sky130_fd_pr__pfet_20v0__tmax_vds_2' SKY130_FD_PR__PFET_20V0__TMAX_VGS_1='100.001n' 
+ SKY130_FD_PR__PFET_20V0__TMAX_VGS_2='20.001n' SKY130_FD_PR__PFET_20V0__VBD_MAX='sky130_fd_pr__pfet_20v0__vbs_max - sky130_fd_pr__pfet_20v0__vds_min' 
+ SKY130_FD_PR__PFET_20V0__VBD_MAX_1='sky130_fd_pr__pfet_20v0__vbs_max - sky130_fd_pr__pfet_20v0__vds_min_1' 
+ SKY130_FD_PR__PFET_20V0__VBD_MAX_2='sky130_fd_pr__pfet_20v0__vbs_max - sky130_fd_pr__pfet_20v0__vds_min_2' 
+ SKY130_FD_PR__PFET_20V0__VBD_MIN='sky130_fd_pr__pfet_20v0__vbs_min' SKY130_FD_PR__PFET_20V0__VBD_MIN_1='sky130_fd_pr__pfet_20v0__vbs_min' 
+ SKY130_FD_PR__PFET_20V0__VBD_MIN_2='sky130_fd_pr__pfet_20v0__vbs_min' SKY130_FD_PR__PFET_20V0__VBD_REVERSEMAX='5.501' 
+ SKY130_FD_PR__PFET_20V0__VBD_REVERSEMIN='-0.501' SKY130_FD_PR__PFET_20V0__VBS_MAX='2.501' 
+ SKY130_FD_PR__PFET_20V0__VBS_MAX_1='2.501' SKY130_FD_PR__PFET_20V0__VBS_MIN='-0.001' 
+ SKY130_FD_PR__PFET_20V0__VBS_MIN_1='-0.001' SKY130_FD_PR__PFET_20V0__VDS_MAX='0.01' 
+ SKY130_FD_PR__PFET_20V0__VDS_MAX_1='0.01' SKY130_FD_PR__PFET_20V0__VDS_MAX_2='0.01' 
+ SKY130_FD_PR__PFET_20V0__VDS_MIN='-28.001' SKY130_FD_PR__PFET_20V0__VDS_MIN_1='-24.501' 
+ SKY130_FD_PR__PFET_20V0__VDS_MIN_2='-24.501' SKY130_FD_PR__PFET_20V0__VGB_MAX='-1*sky130_fd_pr__pfet_20v0__vgs_min' 
+ SKY130_FD_PR__PFET_20V0__VGB_MAX_1='0 + 1.0' SKY130_FD_PR__PFET_20V0__VGB_MAX_2='0 + 1.0' 
+ SKY130_FD_PR__PFET_20V0__VGB_MIN='sky130_fd_pr__pfet_20v0__vgs_min - sky130_fd_pr__pfet_20v0__vbs_max' 
+ SKY130_FD_PR__PFET_20V0__VGB_MIN_1='sky130_fd_pr__pfet_20v0__vgs_min_1 - sky130_fd_pr__pfet_20v0__vbs_max_1' 
+ SKY130_FD_PR__PFET_20V0__VGB_MIN_2='sky130_fd_pr__pfet_20v0__vgs_min_2 - sky130_fd_pr__pfet_20v0__vbs_max_1' 
+ SKY130_FD_PR__PFET_20V0__VGD_MAX='-1*sky130_fd_pr__pfet_20v0__vds_min' SKY130_FD_PR__PFET_20V0__VGD_MAX_1='-1*sky130_fd_pr__pfet_20v0__vds_min_1' 
+ SKY130_FD_PR__PFET_20V0__VGD_MAX_2='-1*sky130_fd_pr__pfet_20v0__vds_min_2' SKY130_FD_PR__PFET_20V0__VGD_MIN='sky130_fd_pr__pfet_20v0__vgs_min' 
+ SKY130_FD_PR__PFET_20V0__VGD_MIN_1='sky130_fd_pr__pfet_20v0__vgs_min_1' SKY130_FD_PR__PFET_20V0__VGD_MIN_2='sky130_fd_pr__pfet_20v0__vgs_min_2' 
+ SKY130_FD_PR__PFET_20V0__VGD_REVERSEMAX='5.501' SKY130_FD_PR__PFET_20V0__VGD_REVERSEMAX_1='0.101' 
+ SKY130_FD_PR__PFET_20V0__VGD_REVERSEMIN='-5.501' SKY130_FD_PR__PFET_20V0__VGD_REVERSEMIN_1='-0.101' 
+ SKY130_FD_PR__PFET_20V0__VGS_MAX='-1*-6.501' SKY130_FD_PR__PFET_20V0__VGS_MAX_1='-1*-5.751' 
+ SKY130_FD_PR__PFET_20V0__VGS_MAX_2='-1*-6.001' SKY130_FD_PR__PFET_20V0__VGS_MIN='-6.501' 
+ SKY130_FD_PR__PFET_20V0__VGS_MIN_1='-5.751' SKY130_FD_PR__PFET_20V0__VGS_MIN_2='-6.001' 
+ SKY130_FD_PR__PFET_20V0__VSD_REVERSEMAX='0.501' SKY130_FD_PR__PFET_20V0__VSD_REVERSEMIN='-5.501' 
+ SKY130_FD_PR__PFET_20V0__VTX='-0.873'
