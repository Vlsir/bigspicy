** Translated using xdm 2.6.0 on Nov_14_2022_16_05_08_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* statistics {
* 	mismatch {
*     	}
*         process {
* 		vary sky130_fd_pr__res_xhigh_po__var_mult dist=gauss std=0.025
* 		vary sky130_fd_pr__res_high_po__var       dist=gauss std=0.025
*         }
* }
.SUBCKT sky130_fd_pr__res_high_po_1p41 r0 r1 b
* .param  w = 1.410 l = 5 mult = 1.0   body_pelgrom = 0.0354   rend_mm = 0.033   rcon = 254.77   rsheet = 230.05   tc1_voltco = -4.68e-3   vc1_body = -1.24e-4   vc2_body = 2.41e-4   vc1_raw_end = -7.62e-2   vc2_raw_end = 0.198   vc3_raw_end = 8.81e-2   r0_var = 15.43   r1_var = 6.96   vc1_end = {vc1_raw_end*0.705/l*(1+tc1_voltco*(temper-30))}   vc2_end = {vc2_raw_end*0.705/l*(1+tc1_voltco*(temper-30))}   vc3_end = {vc3_raw_end*0.705/l*(1+tc1_voltco*(temper-30))}   rtot_var = {sky130_fd_pr__res_high_po__var_mult*sqrt(2*pow(r0_var,2)+pow((r1_var*l),2))}   rend_var = {sky130_fd_pr__res_high_po__var_mult*sqrt(2)*r0_var}   rbody_var = {rtot_var-rend_var}   res_match = {(body_pelgrom/sqrt(w*l*mult))*sky130_fd_pr__res_high_po__slope_spectre}   rend = {(rcon+rend_var)*(1+rend_mm/sqrt(mult)*sky130_fd_pr__res_high_po__con_slope_spectre)}   rbody = {(l*rsheet+rbody_var)*(1+res_match)}; HSpice Parser Retained (as a comment). Continuing.

* rend r0 ra r = {rend*(1+min((abs(v(r0,r1))-1.4),0.6)*vc1_end+pow(min(abs(v(r0,r1))-1.4,0.6),2)*vc2_end+pow(min(abs(v(r0,r1))-1.4,0.6),3)*vc3_end)}; HSpice Parser Retained (as a comment). Continuing.






















* rhrpoly_1p41 ra r1 r = {rbody*(1+abs(v(r0,r1))*vc1_body+pow(abs(v(r0,r1)),2)*vc2_body)}  tc1 = 0.514e-3   tc2 = 0.122e-5; HSpice Parser Retained (as a comment). Continuing.
*+ tnom=30


* c1 r0 b c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_4_1*1e-6)/2}; HSpice Parser Retained (as a comment). Continuing.
* c2 r1 b c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_4_1*1e-6)/2}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__res_high_po_1p41
