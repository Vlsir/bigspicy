** Translated using xdm 2.6.0 on Nov_14_2022_16_05_03_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_MULT=1.0365 SKY130_FD_PR__NFET_05V0_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_05V0_NVT__OVERLAP_MULT=1.1614 SKY130_FD_PR__NFET_05V0_NVT__AJUNCTION_MULT=1.2643e+0 
+ SKY130_FD_PR__NFET_05V0_NVT__PJUNCTION_MULT=1.1856e+0 SKY130_FD_PR__NFET_05V0_NVT__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__WINT_DIFF=2.252e-8 SKY130_FD_PR__NFET_05V0_NVT__DLC_DIFF=-3.0000e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__DWC_DIFF=2.252e-8 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_0=-0.032984 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_0=0.057763 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_0=7.2807e-5 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_0=-0.0067973 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_0=-2.376e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_0=0.021482 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_0=0.0047929 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_0=-1.1063e-18 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_1=-1.119e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_1=0.077833 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_1=0.027909 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_1=-0.002922 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_1=-0.0064693 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_1=-2.2842e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_1=0.013709 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_1=0.0032394 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_2=-1.0808e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_2=-0.14696 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_2=0.0022692 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_2=-0.0072977 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_2=-2.3876e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_2=864.93 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_2=0.027939 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_3=-1.1915e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_3=0.0166 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_3=-8.2319e-19 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_3=0.11551 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_3=0.00089555 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_3=-0.0041127 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_3=-0.0071709 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_3=-0.0033311 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_4=-0.0078839 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_4=0.0084729 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_4=-2.0087e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_4=0.014055 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_4=-1.1143e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_4=0.10719 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_4=0.06314 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_4=-0.0012356 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_5=0.00058708 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_5=-0.0088249 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_5=0.0067298 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_5=-1.6502e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_5=0.019503 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_5=-1.075e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_5=0.11267 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_5=0.088664 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_6=0.044119 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_6=-0.0019442 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_6=-0.0072188 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_6=0.00092262 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_6=-1.3916e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_6=0.0087222 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_6=-9.064e-19 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_6=0.13457 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_7=-0.032084 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_7=0.00069292 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_7=-0.0092302 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_7=0.0096456 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_7=-1.9874e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_7=288.71 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_7=-1.0787e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_8=0.041165 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_8=4.35e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_8=0.00055638 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_8=-0.010837 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_8=-0.010299 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_8=-2.8046e-12 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_8=3.3176e-10 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_8=-7.4006e-19 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_9=0.13133 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_9=0.0023042 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_9=-0.01127 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_9=0.020187 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_9=4.2431e-12 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_9=-4479.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_9=-3.7969e-19 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_10=-1768.2 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_10=0.013913 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_10=0.0061791 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_10=-0.010406 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_10=0.00086128 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_10=-1.3004e-11 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_10=-8.7248e-19 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0, L = 2.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0, L = 4.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0, L = 0.9
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0, L = 25.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0, L = 2.0
* ------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0, L = 4.0
* ------------------------------------
*














* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0, L = 8.0
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0, L = 0.9
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42, L = 1.0
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42, L = 0.9
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7, L = 0.9
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_05v0_nvt.pm3.spice




















