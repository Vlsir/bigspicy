** Translated using xdm 2.6.0 on Nov_14_2022_16_05_31_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PFET_01V8__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__pfet_01v8 d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__pfet_01v8 d g s b sky130_fd_pr__pfet_01v8__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__pfet_01v8__model.0 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.069382+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43448553   k2 = 0.018008346   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.6113816e-10   ub = 7.7273446e-19   uc = -6.6549964e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0097753   a0 = 1.33379   keta = 0.0051290095   a1 = 0.0   a2 = 0.9995   ags = 0.1474578   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22144045+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.2879038+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0015228006   pdiblc1 = 0.39   pdiblc2 = 0.0029632464   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.3760948e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.6464006   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1181082000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4485   kt2 = -0.0075706   at = 90900.0   ute = -0.33954   ua1 = 1.6104e-9   ub1 = -5.609e-19   uc1 = -1.0858e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.1 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.069382+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43448553   k2 = 0.018008346   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.6113816e-10   ub = 7.7273446e-19   uc = -6.6549964e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0097753   a0 = 1.33379   keta = 0.0051290095   a1 = 0.0   a2 = 0.9995   ags = 0.1474578   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22144045+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.2879038+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0015228006   pdiblc1 = 0.39   pdiblc2 = 0.0029632464   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.3760948e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.6464006   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1181082000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4485   kt2 = -0.0075706   at = 90900.0   ute = -0.33954   ua1 = 1.6104e-9   ub1 = -5.609e-19   uc1 = -1.0858e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.2 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.071713954212+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.88017026439316e-8   k1 = 0.438164888574485 lk1 = -2.96653362582688e-8   k2 = 0.016478384967666 lk2 = 1.23355219578153e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 268861.1090625 lvsat = -0.875188140274457   ua = -5.7232489780447e-10 lua = 9.01946173183564e-17   ub = 7.87456738993755e-19 lub = -1.18700406061651e-25   uc = -7.3282823639794e-11 luc = 5.42846099804694e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0096601242127 lu0 = 9.28620679364886e-10   a0 = 1.474672129245 la0 = -1.13588160877165e-6   keta = 0.0215972828408877 lketa = -1.32777726432629e-07 pketa = 1.0097419586829e-28   a1 = 0.0   a2 = 1.20212407025 la2 = -1.63368452851232e-6   ags = 0.0341385976396201 lags = 9.1365170708049e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.227497548716745+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.88361942833796e-8   nfactor = {1.11405915264415+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.40164645986788e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.437343739836769 lpclm = 3.53842204585403e-06 wpclm = -3.63959469523332e-23 ppclm = -3.66031460022549e-28   pdiblc1 = 0.39   pdiblc2 = 0.00581349077122623 lpdiblc2 = -2.29804885767347e-8   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.01483080305984e-08 lpscbe2 = -6.22607573712542e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.2324138664649 lbeta0 = 1.1400463169296e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 8.4131752392395e-11 lagidl = 1.27939936154485e-16   bgidl = 1364999653.579 lbgidl = -1482.86146261688   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.43142804353597 lkt1 = -1.37645004921234e-7   kt2 = 0.00995327517421449 lkt2 = -1.41288661886878e-7   at = 87833.957571185 lat = 0.0247203901961761   ute = -0.47558397427718 lute = 1.09687331667821e-6   ua1 = 1.22054489018415e-09 lua1 = 3.14326062289545e-15   ub1 = -2.9714671580816e-19 lub1 = -2.12654725174993e-24   uc1 = -8.812855842886e-11 luc1 = -1.64892569966253e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.3 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0736386915303+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.66212136132752e-8   k1 = 0.42415958432975 lk1 = 2.72331449679531e-8   k2 = 0.021881869435854 lk2 = -9.61687937505504e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53437.5   ua = -2.2098226734349e-10 lua = -1.33718330421238e-15   ub = 5.0506631000493e-19 lub = 1.02854968158465e-24   uc = -8.1250014202858e-11 luc = 8.66524211152146e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01110981263557 lu0 = -4.96093859554684e-9   a0 = 1.215236098536 la0 = -8.18869318440973e-8   keta = -0.00536872903134401 lketa = -2.32245818920487e-8   a1 = 0.0   a2 = 0.8   ags = 0.0616891254330901 lags = 8.01723885946682e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22143888795771+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.4222048854615e-8   nfactor = {1.4671344584266+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.27706942655251e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.1619898605 leta0 = -3.33095122881999e-7   etab = -0.141676670056533 letab = 2.91196363485133e-7   dsub = 0.8693957 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = 0.46514143279979 lpclm = -1.28048510935813e-7   pdiblc1 = 0.39   pdiblc2 = -2.46391392811899e-05 lpdiblc2 = 7.37719846629315e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800453914.43147 lpscbe1 = -1.84409001803806   pscbe2 = 8.2808066288523e-09 lpscbe2 = 1.36090642266155e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.8583712272946 lbeta0 = 8.85742500880952e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.3173649521521e-10 lagidl = -6.54609010177104e-17 wagidl = 1.97215226305253e-31   bgidl = 915838594.2136 lbgidl = 341.917325281249   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.46638552985471 lkt1 = 4.37460738175925e-9   kt2 = -0.00514777539406101 lkt2 = -7.99385600082808e-8   at = 107262.402188066 lat = -0.0542103471852601   ute = -0.17519952681143 lute = -1.23479954205146e-7   ua1 = 2.3512472320185e-09 lua1 = -1.45037367772978e-15   ub1 = -1.03511635614758e-18 lub1 = 8.71556251939332e-25   uc1 = -2.44462937652451e-10 luc1 = 4.70237419773918e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.4 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0810491947134+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.19063990778584e-8   k1 = 0.3517509538705 lk1 = 1.7658593768116e-7   k2 = 0.050734812238536 lk2 = -6.91300556116934e-08 pk2 = 5.04870979341448e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 34509.260625 lvsat = 0.0390421058079712   ua = -7.41991490889919e-10 lua = -2.62529881375017e-16   ub = 9.5358754654408e-19 lub = 1.03412735292012e-25   uc = -4.311338214219e-11 luc = 7.99035463486248e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00938543840832 lu0 = -1.40417878820035e-9   a0 = 1.339169500344 la0 = -3.37516675882548e-7   keta = -0.00634552755000199 lketa = -2.1209800149121e-8   a1 = 0.0   a2 = 0.6937362 la2 = 2.191837519044e-7   ags = 0.3200841249827 lags = 2.68748540865674e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.2244805575492+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.04959121374668e-8   nfactor = {1.1842794114134+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.50656874195687e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.519661301 leta0 = 1.07290446557204e-06 weta0 = 1.15805285757424e-23 peta0 = 3.47098798297245e-28   etab = 7.90303547058587 letab = -1.63021325968652e-05 wetab = 1.07698915754404e-21 petab = -8.10160149661979e-27   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = 0.17517350209466 lpclm = 4.70050361717955e-7   pdiblc1 = 0.40922897655538 lpdiblc1 = -3.9662417744236e-8   pdiblc2 = 0.00022996388166064 lpdiblc2 = 2.12565980719901e-10   pdiblcb = -0.0507746564432779 lpdiblcb = 5.31637858168499e-8   drout = 0.39466727773572 ldrout = 3.4102155558575e-7   pscbe1 = 799092171.13706 lpscbe1 = 0.964693447256877   pscbe2 = 8.9459879377396e-09 lpscbe2 = -1.1121821939135e-17   pvag = 0.0   delta = 0.01   alpha0 = -4.7443750631206e-05 lalpha0 = 9.78594891782495e-11 walpha0 = 7.17685930047446e-27 palpha0 = 2.04423169585399e-32   alpha1 = 2.062638e-10 lalpha1 = -2.191837519044e-16   beta0 = -14.951711701752 lbeta0 = 4.76558168414124e-05 pbeta0 = -2.58493941422821e-26   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 788249290.6404 lbgidl = 605.087871224867   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.45593337680516 lkt1 = -1.71844006800584e-8   kt2 = -0.040229346696406 lkt2 = -7.57797794035452e-9   at = 70516.470352408 lat = 0.0215832081643779   ute = -0.16229860395988 lute = -1.50089887913821e-7   ua1 = 1.4080917459452e-09 lua1 = 4.95014667753484e-16   ub1 = 1.13857555640005e-20 lub1 = -1.28699877075722e-24   uc1 = -2.1779306702286e-11 luc1 = 1.09217005981318e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.5 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0806963110872+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.15314115270799e-8   k1 = 0.56579981919688 lk1 = -5.08705204715343e-8   k2 = -0.035713367390328 lk2 = 2.27330650927634e-08 wk2 = 2.64697796016969e-23   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 61674.84647184 lvsat = 0.0101749219948569   ua = -6.15372854171e-10 lua = -3.97079656260737e-16   ub = 8.2648775408584e-19 lub = 2.38473804550251e-25   uc = -6.0901074890088e-11 luc = 2.68922328811033e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00945805566708 lu0 = -1.48134464681456e-9   a0 = 1.147070287248 la0 = -1.3338475227664e-7   keta = -0.0444291047069 lketa = 1.92592561137308e-8   a1 = 0.0   a2 = 1.0125276 la2 = -1.195761038088e-7   ags = 0.27373978293884 lags = 3.17995799806477e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.18356061611124+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.29871725922842e-8   nfactor = {1.7660613454352+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.75667166093699e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -15.8080632511956 letab = 8.89418192665119e-6   dsub = 0.21572307880964 ldsub = 4.70503389798817e-8   voffl = 0.0   minv = 0.0   pclm = 0.61122775131572 lpclm = 6.68254643418589e-9   pdiblc1 = 0.746679578145028 lpdiblc1 = -3.98250250116256e-7   pdiblc2 = 0.00043   pdiblcb = 0.251604512886556 lpdiblcb = -2.68155809921466e-07 wpdiblcb = -1.32348898008484e-23 ppdiblcb = 7.65195078064381e-29   drout = 0.39554400452856 ldrout = 3.4008991238006e-7   pscbe1 = 800000000.0   pscbe2 = 8.6986084540396e-09 lpscbe2 = 2.5175301786087e-16   pvag = 0.0   delta = 0.01   alpha0 = 9.4887801262412e-05 lalpha0 = -5.3387426462881e-11   alpha1 = -1.125276e-10 lalpha1 = 1.195761038088e-16   beta0 = 52.9527565495392 lbeta0 = -2.45020514922032e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1741875147.7596 lbgidl = -408.271202332566   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.43119522972308 lkt1 = -4.34720958190658e-8   kt2 = -0.03855268902226 lkt2 = -9.35965809789368e-9   at = 108637.67837344 lat = -0.0189258360846755   ute = -0.22847566465708 lute = -7.97676284886699e-8   ua1 = 3.4706461072424e-09 lua1 = -1.69673397362665e-15   ub1 = -3.0145161509524e-18 lub1 = 1.92843957937956e-24   uc1 = -5.1810348954744e-11 luc1 = 4.28338272751993e-17 wuc1 = 2.46519032881566e-32 puc1 = -2.35098870164458e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.6 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0341750978416+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.53568091490022e-8   k1 = 0.03869703848784 lk1 = 2.45697533861039e-7   k2 = 0.15332470314536 lk2 = -8.3626936837295e-08 wk2 = 1.05879118406788e-22 pk2 = -4.41762106923767e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93447.90228032 lvsat = -0.00770180657911469   ua = -4.781111169976e-10 lua = -4.74308325540504e-16   ub = 4.01574301748799e-19 lub = 4.77546259546259e-25   uc = -2.96125602439574e-11 luc = 9.28812557763372e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0094312253128 lu0 = -1.46624886994317e-9   a0 = 1.22837436956264 la0 = -1.79129518541985e-07 wa0 = -1.6940658945086e-21   keta = 0.079523086206992 lketa = -5.04809566776795e-08 wketa = 5.29395592033938e-23   a1 = 0.0   a2 = 0.8   ags = -0.67367344200792 lags = 8.51046481864072e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20928156205992+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.48440899438927e-9   nfactor = {0.8301648484944+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 4.59004216636408e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.10067225483276 leta0 = -3.43587416114595e-7   etab = 0.0061540160017152 letab = -3.49764813017304e-09 wetab = -6.20385459414771e-25 petab = 2.95822839457879e-31   dsub = 0.1527052563208 ldsub = 8.25065605893578e-8   voffl = 0.0   minv = 0.0   pclm = 0.43613961756656 lpclm = 1.05193783830546e-7   pdiblc1 = -0.440678271693176 lpdiblc1 = 2.69802395801011e-07 ppdiblc1 = -1.0097419586829e-28   pdiblc2 = -0.011651542854336 lpdiblc2 = 6.7975351084779e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = 2.76101316827354e-30   pdiblcb = -0.4125828 lpdiblcb = 1.055412114264e-7   drout = 1.66428035421992 ldrout = -3.73749369937587e-7   pscbe1 = 800004426.95408 lpscbe1 = -0.002490772589681   pscbe2 = 9.47692126902e-09 lpscbe2 = -1.86155347734076e-16   pvag = 0.0   delta = 0.01   alpha0 = -9.95210267414e-09 lalpha0 = 5.65569494437278e-15 walpha0 = 1.38050658413677e-30 palpha0 = 2.53906779777614e-36   alpha1 = 2.250552e-10 lalpha1 = -7.03608076176e-17   beta0 = 1.6659968511696 lbeta0 = 4.35382841096804e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 333261981.0512 lbgidl = 384.268092557915   cgidl = 592.646478140784 lcgidl = -0.000164654029168174   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.44538215712 lkt1 = -3.54899913623174e-8   kt2 = 0.028313858144 lkt2 = -4.69813184624239e-8   at = 59993.376 lat = 0.008443296914112   ute = -0.379316502 lute = 5.10115855227605e-9   ua1 = 8.555843332e-10 lua1 = -2.25400847202982e-16   ub1 = 4.3834119456e-19 lub1 = -1.42691717848492e-26   uc1 = 7.23120692000001e-12 luc1 = 9.61480436094503e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.7 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.990413833542857+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.67537500117172e-9   k1 = 0.139611906368572 lk1 = 2.14147711396542e-7   k2 = 0.139717634085772 lk2 = -7.93728499806434e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 13145.6035371429 lvsat = 0.0174037434953547   ua = -1.07630223388571e-09 lua = -2.87291051138838e-16   ub = 1.01120439936571e-18 lub = 2.86952725087502e-25   uc = -1.07347336365771e-13 luc = 6.3674824630078e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00674226626085715 lu0 = -6.25578089861856e-10   a0 = 1.08482302099057 la0 = -1.3424991202711e-7   keta = -0.284954641152943 lketa = 6.34686310486757e-8   a1 = 0.0   a2 = 0.898081940028286 la2 = -3.06641415665632e-8   ags = 4.81618663288 lags = -8.65292392228738e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0589799012225715+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.55056016464777e-8   nfactor = {4.07603463828571+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -5.55778022704369e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.584620529535577 leta0 = 1.83299149404753e-07 weta0 = -7.27918939046664e-23 peta0 = 8.83524213847533e-29   etab = 0.175871445820531 letab = -5.65577659538681e-08 petab = -1.26217744835362e-29   dsub = 0.879662738218 ldsub = -1.44767972636019e-7   voffl = 0.0   minv = 0.0   pclm = 1.24484513952457 lpclm = -1.47638293143363e-7   pdiblc1 = 1.23931561133057 lpdiblc1 = -2.55427531799767e-7   pdiblc2 = 0.0306017834527886 lpdiblc2 = -6.41246032152891e-9   pdiblcb = -0.075   drout = -1.19818899299457 ldrout = 5.21167321836857e-7   pscbe1 = 799984189.449715 lpscbe1 = 0.00383624030018836   pscbe2 = 7.77486197647142e-09 lpscbe2 = 3.45973065369725e-16   pvag = 0.0   delta = 0.01   alpha0 = 3.60003666933571e-08 lalpha0 = -8.71079317374279e-15   alpha1 = -3.46625714285714e-10 lalpha1 = 1.08368370062857e-16   beta0 = 39.81024323392 lbeta0 = -7.57151248964228e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.49192114402857e-11 lagidl = 1.4093967573732e-17   bgidl = 3511720739.85429 lbgidl = -609.438896876764   cgidl = -745.165993359943 lcgidl = 0.00025359698629687 wcgidl = -4.33680868994202e-19   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.5589   kt2 = -0.12196   at = 256846.6 lat = -0.0531005013308   ute = -0.5813742 lute = 6.82720731396e-8   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 3.7985e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.8 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.932957859466665+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.22656276367267e-8   k1 = -0.86434125910667 lk1 = 4.57744899561124e-7   k2 = 0.570090003164 lk2 = -1.83797540869047e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 294060.394053333 lvsat = -0.0507568594459127   ua = -6.46665128013335e-10 lua = -3.91537339233501e-16   ub = 7.44576124093334e-19 lub = 3.51646876543041e-25   uc = 3.25316059937333e-13 luc = -4.13057565221147e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00808365713333333 lu0 = -9.51050488377733e-10   a0 = -1.430645407812 la0 = 4.76098316600688e-7   keta = -0.124531741410173 lketa = 2.45439395008896e-8   a1 = 0.0   a2 = -0.842900560066002 la2 = 3.91764370291314e-7   ags = 1.25   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0908657602386662+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.77688805865304e-8   nfactor = {1.750172092+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 8.56461380130426e-9   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.998252372324667 leta0 = 2.83661952475413e-7   etab = -0.338688758357333 letab = 6.82940928674407e-08 wetab = -4.2351647362715e-22 petab = 1.0097419586829e-28   dsub = 0.446191827990666 ldsub = -3.95914579202794e-8   voffl = 0.0   minv = 0.0   pclm = 2.83441603732867 lpclm = -5.33328596644753e-7   pdiblc1 = 1.37103628340867 lpdiblc1 = -2.87387972231452e-7   pdiblc2 = 0.0307086957296267 lpdiblc2 = -6.43840130255636e-09 ppdiblc2 = 6.31088724176809e-30   pdiblcb = -0.584736382052253 lpdiblcb = 1.23681416268395e-7   drout = 0.593438031821332 ldrout = 8.64505237895754e-8   pscbe1 = 899843393.227332 lpscbe1 = -24.2258012458938   pscbe2 = 1.058390275688e-08 lpscbe2 = -3.35606971507051e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 17.3103286992 lbeta0 = -2.11217822676689e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.05188506639333e-10 lagidl = -2.23670736747746e-17   bgidl = 675055822.713332 lbgidl = 78.8438052884821   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.370328060000001 lkt1 = -2.2546603802228e-7   kt2 = -0.12196   at = 38000.0   ute = -0.3   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 3.7985e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.9 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.07842466109461+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.25846390360971e-8   k1 = 0.444135669148989 wk1 = -6.6789020286023e-8   k2 = 0.0135611189666637 wk2 = 3.07794459707013e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.84872715608765e-10 wua = 1.64267860966509e-16   ub = 8.63568902318425e-19 wub = -6.28669008499281e-25   uc = -7.47240562252678e-11 wuc = 5.65732372377703e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.010383319369021 wu0 = -4.20812771141171e-9   a0 = 1.557033079403 wa0 = -1.54507477340611e-6   keta = 0.0297110219689129 wketa = -1.70133145658272e-7   a1 = 0.0   a2 = 1.22027301148113 wa2 = -1.527979329082e-6   ags = 0.047081358434931 wags = 6.94709587957677e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.230934813558148+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 6.57108908480845e-8   nfactor = {0.71646106133894+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.95497930915677e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.5539667051391 wpclm = 3.84456631087745e-6   pdiblc1 = 0.39   pdiblc2 = 0.00983928660989256 wpdiblc2 = -4.75893644615633e-8   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.01118663929499e-08 wpscbe2 = -5.09230624436736e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 0.451794529844371 wbeta0 = 2.90310456239233e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 292047992.46066 wbgidl = 6153.04188341489   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.479124531398196 wkt1 = 2.11953674162139e-7   kt2 = 0.0981458514558926 wkt2 = -7.31668021760484e-7   at = 93114.46899 wat = -0.0153264333303815   ute = -0.769707712213479 wute = 2.97720888930694e-6   ua1 = 7.51784184559411e-10 wua1 = 5.94251629225174e-15   ub1 = -8.96433815969241e-20 wub1 = -3.26158694299698e-24   uc1 = -6.51151131704926e-10 wuc1 = 3.75515769903155e-15   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.10 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.07842466109461+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.25846390360971e-8   k1 = 0.444135669148989 wk1 = -6.67890202860247e-8   k2 = 0.0135611189666637 wk2 = 3.07794459707013e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 160312.5   ua = -5.84872715608765e-10 wua = 1.6426786096651e-16   ub = 8.63568902318425e-19 wub = -6.28669008499287e-25   uc = -7.47240562252678e-11 wuc = 5.65732372377703e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.010383319369021 wu0 = -4.20812771141174e-9   a0 = 1.557033079403 wa0 = -1.54507477340611e-6   keta = 0.0297110219689129 wketa = -1.70133145658272e-7   a1 = 0.0   a2 = 1.22027301148113 wa2 = -1.527979329082e-6   ags = 0.0470813584349311 wags = 6.94709587957677e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.230934813558148+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 6.57108908480845e-8   nfactor = {0.716461061338941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.95497930915677e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.553966705139099 wpclm = 3.84456631087745e-6   pdiblc1 = 0.39   pdiblc2 = 0.00983928660989256 wpdiblc2 = -4.75893644615633e-8   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.01118663929499e-08 wpscbe2 = -5.09230624436731e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 0.451794529844367 wbeta0 = 2.90310456239233e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 292047992.46066 wbgidl = 6153.04188341489   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.479124531398196 wkt1 = 2.11953674162139e-7   kt2 = 0.0981458514558926 wkt2 = -7.31668021760484e-7   at = 93114.46899 wat = -0.0153264333303813   ute = -0.769707712213479 wute = 2.97720888930694e-6   ua1 = 7.51784184559411e-10 wua1 = 5.94251629225174e-15   ub1 = -8.96433815969241e-20 wub1 = -3.26158694299699e-24   uc1 = -6.51151131704926e-10 wuc1 = 3.75515769903155e-15   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.11 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08189368379834+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.7969474273919e-08 wvth0 = 7.04543380516281e-08 pvth0 = -6.34505343311321e-14   k1 = 0.417809114724208 lk1 = 2.12261478114308e-07 wk1 = 1.40883169831425e-07 pk1 = -1.67438569158417e-12   k2 = 0.0208387755148587 lk2 = -5.86771102364261e-08 wk2 = -3.01784469856019e-08 pk2 = 4.91481424149423e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 277173.547059667 lvsat = -0.942208318743057 wvsat = -0.057530734163274 pvsat = 4.63849483432709e-7   ua = -2.36391719402569e-10 lua = -2.80967612228993e-15 wua = -2.32500770409969e-15 pua = 2.00701277633742e-20   ub = 7.06167150986329e-19 lub = 1.26907334155671e-24 wub = 5.62608669020016e-25 pub = -9.60484067131883e-30   uc = -9.29444964213673e-11 luc = 1.46904813501799e-16 wuc = 1.3607926704386e-16 puc = -6.41028337143709e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0119721469262656 lu0 = -1.28101414384876e-08 wu0 = -1.60016067679461e-08 pu0 = 9.50865523934186e-14   a0 = 2.00018050141977 la0 = -3.57293724435446e-06 wa0 = -3.63706562027491e-06 pa0 = 1.68669648976165e-11   keta = 0.0727536623029575 lketa = -3.47037227577601e-07 wketa = -3.54055461056198e-07 pketa = 1.4828990491753e-12   a1 = 0.0   a2 = 1.64712728818555 la2 = -3.44157151181958e-06 wa2 = -3.07988605046776e-06 pa2 = 1.25124621043002e-11   ags = -0.133360671356584 lags = 1.4548387661942e-06 wags = 1.15926950919188e-06 pags = -3.74557847421991e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.254443439561762+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.89541541344528e-07 wvoff = 1.86493647654957e-07 pvoff = -9.73827644775852e-13   nfactor = {0.132709470345201+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.70657776010657e-06 wnfactor = 6.79196256414761e-06 pnfactor = -2.28735689970529e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.54053419600524 lpclm = 7.95433654142196e-06 wpclm = 7.63522770177921e-06 ppclm = -3.05627305754173e-11   pdiblc1 = 0.39   pdiblc2 = 0.0195496752619774 lpdiblc2 = -7.82913485410683e-08 wpdiblc2 = -9.50687125274746e-08 ppdiblc2 = 3.82808795931443e-13   pdiblcb = -0.025   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.37544635861039e-08 lpscbe2 = -2.93689425482167e-14 wpscbe2 = -2.49583547794178e-14 ppscbe2 = 1.60172757828542e-19   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -3.64445705592367 lbeta0 = 3.30265936929736e-05 wbeta0 = 4.75951138578042e-05 pbeta0 = -1.49675361977081e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.50875943338585e-11 lagidl = 4.42738848595249e-16 wagidl = 2.70226265586602e-16 pagidl = -2.17873655751663e-21   bgidl = 789132801.642863 lbgidl = -4007.81487173519 wbgidl = 3985.59878383115 pbgidl = 0.0174753090975417   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.487056361199977 lkt1 = 6.39514723693706e-08 wkt1 = 3.85005934067596e-07 pkt1 = -1.3952577266996e-12   kt2 = 0.156558599634276 lkt2 = -4.70960843147468e-07 wkt2 = -1.01466163733278e-06 pkt2 = 2.28167507867059e-12   at = 93304.5908732254 lat = -0.00153288392032414 wat = -0.0378624839441466 pat = 1.81700018048467e-7   ute = -1.34264958727912 lute = 4.61942293369546e-06 wute = 6.00099769775527e-06 pute = -2.43797145509702e-11   ua1 = -4.25639234427394e-11 lua1 = 6.40454124080623e-15 wua1 = 8.74202940230362e-15 pua1 = -2.25714607826026e-20   ub1 = 3.96333870400639e-19 lub1 = -3.91825865909113e-24 wub1 = -4.79960840203184e-24 pub1 = 1.24005102604299e-29   uc1 = -1.18582959783409e-09 luc1 = 4.31091891879473e-15 wuc1 = 7.59723521670748e-15 puc1 = -3.09772801929596e-20   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.12 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0786304006128+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.47119359995876e-08 wvth0 = 3.45478292100828e-08 pvth0 = 8.24246129358626e-14   k1 = 0.515358872049934 lk1 = -1.84047872887965e-07 wk1 = -6.31194118921337e-07 pk1 = 1.46228484063977e-12   k2 = -0.0112270279384703 lk2 = 7.15946413735995e-08 wk2 = 2.29148075923168e-07 pk2 = -5.62068362227614e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 36812.6240056666 lvsat = 0.0342911009711996 wvsat = 0.115061468326548 pvsat = -2.37330156906133e-7   ua = -1.27890995349834e-09 lua = 1.42569807124043e-15 wua = 7.32196216042606e-15 pua = -1.91220185931029e-20   ub = 1.25066766677043e-18 lub = -9.43035144887378e-25 wub = -5.16033845455129e-24 pub = 1.36454217848926e-29   uc = -6.26323506940766e-11 luc = 2.37575384085707e-17 wuc = -1.28853634809675e-16 puc = 4.35298137376732e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00752896053312475 lu0 = 5.24091644336942e-09 wu0 = 2.47832285129823e-08 pu0 = -7.0607469242622e-14   a0 = 1.07594511511541 la0 = 1.81896556990304e-07 wa0 = 9.6403877433338e-07 pa0 = -1.82565665788613e-12   keta = -0.00888046890715201 lketa = -1.53873040264241e-08 wketa = 2.43048998758902e-08 pketa = -5.4242130841114e-14   a1 = 0.0   a2 = 0.8   ags = -0.0380112822827168 lags = 1.06746871486592e-06 wags = 6.90030729158303e-07 pags = -1.83923117538186e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.213699127766288+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.40121519603848e-08 wvoff = -5.3567206902714e-08 pvoff = 1.45270526261525e-15   nfactor = {0.781719525969132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.06988484574666e-06 wnfactor = 4.74378567204827e-06 pnfactor = -1.45525677244882e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.161989865346782 leta0 = -3.33095142572719e-07 weta0 = -3.35447823828655e-14 peta0 = 1.36280307321984e-19   etab = -0.141676670031157 letab = 2.9119636338204e-07 wetab = -1.75627199415496e-16 petab = 7.13509517399476e-22   dsub = 0.869395700000001 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = 1.03107602397316 lpclm = -2.49318485945064e-06 wpclm = -3.91685718795067e-06 ppclm = 1.6369208476825e-11   pdiblc1 = 0.39   pdiblc2 = 0.000468599967088319 lpdiblc2 = -7.71846967190569e-10 wpdiblc2 = -3.41372866987366e-09 ppdiblc2 = 1.0447775622167e-14   pdiblcb = -0.025   drout = 0.56   pscbe1 = 772264117.218925 lpscbe1 = 112.680851349933 wpscbe1 = 195.102776117452 ppscbe1 = -0.000792631952160262   pscbe2 = 5.33982481412947e-09 lpscbe2 = 4.8166886830798e-15 wpscbe2 = 2.03546592491293e-14 ppscbe2 = -2.39176148583661e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 0.905519129316168 lbeta0 = 1.45416875437232e-05 wbeta0 = 2.04368139804672e-05 pbeta0 = -3.93410208800167e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.09824811332283e-10 lagidl = -2.26528829196798e-16 wagidl = -5.40452531173204e-16 pagidl = 1.11475792799404e-21   bgidl = -847450994.08005 lbgidl = 2641.03264695295 wbgidl = 12203.801651401 pbgidl = -0.0159122741639564   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.481191257039958 lkt1 = 4.01236773349203e-08 wkt1 = 1.0247106265079e-07 pkt1 = -2.47420821756572e-13   kt2 = 0.125542580920162 lkt2 = -3.44953986910796e-07 wkt2 = -9.04513471183775e-07 pkt2 = 1.83418295324332e-12   at = 101602.825215108 lat = -0.0352456060905637 wat = 0.0391701710639873 pat = -1.31255773428466e-7   ute = -0.32667543599748 lute = 4.91887739680936e-07 wute = 1.04837115976002e-06 pute = -4.25898577790225e-12   ua1 = 1.03899214991823e-09 lua1 = 2.01057043803918e-15 wua1 = 9.08217280038044e-15 pua1 = -2.39533402770786e-20   ub1 = -3.60387251747629e-19 lub1 = -8.43974672848933e-25 wub1 = -4.66982860512026e-24 pub1 = 1.18732619258646e-29   uc1 = 9.49632295322931e-11 luc1 = -8.92478691791384e-16 wuc1 = -2.34918282686987e-15 puc1 = 9.43141571476337e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.13 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.11550155001117+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.076376985235e-08 wvth0 = 2.38446204905273e-07 pvth0 = -3.38143924911313e-13   k1 = 0.321412563560375 lk1 = 2.15993152962322e-07 wk1 = 2.09973279616448e-07 pk1 = -2.72738999945413e-13   k2 = 0.0696936020775574 lk2 = -9.53153250813998e-08 wk2 = -1.31214584536798e-07 pk2 = 1.81229355018209e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -78668.674762849 lvsat = 0.272487216100493 wvsat = 0.783309266928176 pvsat = -1.6156834597182e-6   ua = -5.0840183122702e-10 lua = -1.63581261065036e-16 wua = -1.61668389201057e-15 pua = -6.84827576797165e-22   ub = 8.54356158651336e-19 lub = -1.25587968403626e-25 wub = 6.86784623170246e-25 pub = 1.58492353410721e-30   uc = -5.35724710392645e-11 luc = 5.07028635712815e-18 wuc = 7.2387795630204e-17 puc = 2.02099157770806e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0111556698579779 lu0 = -2.23967202502708e-09 wu0 = -1.22518465668496e-08 pu0 = 5.7824839498924e-15   a0 = 0.590790142439593 la0 = 1.18259563952041e-06 wa0 = 5.1795651176653e-06 pa0 = -1.05207614836436e-11   keta = -0.0734570185504656 lketa = 1.17810741176761e-07 wketa = 4.64481461319129e-07 pketa = -9.62167033183273e-13   a1 = 0.0   a2 = 0.432271877933821 la2 = 7.58489998242341e-07 wa2 = 1.80960560681442e-06 pa2 = -3.73256128962849e-12   ags = 1.80783979922172 lags = -2.73985386818622e-06 wags = -1.02968198046977e-05 pags = 2.08226642360698e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.208872001906996+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.40555387322272e-08 wvoff = -1.08027472280742e-07 pvoff = 1.13784518121421e-13   nfactor = {2.15638577474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.65553996285577e-07 wnfactor = -6.72798916347195e-06 pnfactor = 9.10955097869958e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.519661310693564 leta0 = 1.07290447587279e-06 weta0 = 6.70895648087443e-14 peta0 = -7.12919206757202e-20   etab = 27.3478901066646 letab = -5.64098286737681e-05 wetab = -0.000134578659509167 petab = 2.77587057093019e-10   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = -1.53717203027296 lpclm = 2.80418117066348e-06 wpclm = 1.18512156904978e-05 ppclm = -1.61546178290321e-11   pdiblc1 = 0.433691578527892 lpdiblc1 = -9.01199101516136e-08 wpdiblc1 = -1.69306700573559e-07 ppdiblc1 = 3.49218434257643e-13   pdiblc2 = -0.000262229208275453 lpdiblc2 = 7.3558906142341e-10 wpdiblc2 = 3.40648914599609e-09 ppdiblc2 = -3.619864813123e-15   pdiblcb = -0.0508216502364223 lpdiblcb = 5.32607170003536e-08 wpdiblcb = 3.25246025490097e-10 ppdiblcb = -6.7086481152505e-16   drout = 0.646469185779945 ldrout = -1.78354628418774e-07 wdrout = -1.74273163161459e-06 pdrout = 3.59462448717027e-12   pscbe1 = 855471765.562147 lpscbe1 = -58.9464060134278 wpscbe1 = -390.205552234907 ppscbe1 = 0.0004146472476158   pscbe2 = 1.82363132192383e-09 lpscbe2 = 1.20693229954558e-14 wpscbe2 = 4.92941307015101e-14 ppscbe2 = -8.3609268375962e-20   pvag = 0.0   delta = 0.01   alpha0 = -0.000164180346174537 lalpha0 = 3.38644827136554e-10 walpha0 = 8.07938904039724e-10 palpha0 = -1.66648548515069e-15   alpha1 = 4.6772812206618e-10 lalpha1 = -7.58489998242342e-16 walpha1 = -1.80960560681442e-15 palpha1 = 3.73256128962849e-21   beta0 = -70.1725880342572 lbeta0 = 0.000161150092347382 wbeta0 = 0.00038218601541825 pbeta0 = -7.85498670235242e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = -1005300637.85486 lbgidl = 2966.61932048933 wbgidl = 12413.2347429227 pbgidl = -0.0163442588169865   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.455710751183931 lkt1 = -1.24333823029437e-08 wkt1 = -1.54080131932718e-09 pkt1 = -3.28819986809815e-14   kt2 = -0.036596980431235 lkt2 = -1.05187663640731e-08 wkt2 = -2.51397602071055e-08 pkt2 = 2.03533207818281e-14   at = -93219.77422522 lat = 0.366602890773836 wat = 1.13322545839128 pat = -2.38789578317067e-6   ute = 0.306950422346337 lute = -8.15053033521638e-07 wute = -3.24769231337424e-06 pute = 4.60223799219645e-12   ua1 = 2.24293785270969e-09 lua1 = -4.72733718475201e-16 wua1 = -5.77800513542274e-15 pua1 = 6.69782742007062e-21   ub1 = -4.10626663507795e-19 lub1 = -7.40348953054769e-25 wub1 = 2.92076576131998e-24 pub1 = -3.78338645694097e-30   uc1 = -6.8356343669916e-10 luc1 = 7.13339993990929e-16 wuc1 = 4.58023589099865e-15 puc1 = -4.86146665062353e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.14 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.07256075278565+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.51332469702156e-08 wvth0 = -5.63065423256088e-08 pvth0 = -2.49284550993943e-14   k1 = 0.596985343184793 lk1 = -7.68409544322104e-08 wk1 = -2.15836327549457e-07 pk1 = 1.79742469394154e-13   k2 = -0.0524881483644272 lk2 = 3.45196458447699e-08 wk2 = 1.16098967017498e-07 pk2 = -8.15754227783449e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 283779.388816549 lvsat = -0.112663869285391 wvsat = -1.53719491037942 pvsat = 8.50172458247589e-7   ua = -6.82912452943618e-12 lua = -6.96571478964743e-16 wua = -4.21175683339465e-15 pua = 2.07279554348935e-21   ub = 3.41145619726734e-19 lub = 4.19769052258136e-25 wub = 3.35907339333744e-24 pub = -1.25475206004572e-30   uc = -8.56306944158944e-11 luc = 3.91365727296234e-17 wuc = 1.7115474032805e-16 puc = -8.47435928027493e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0107518121265683 lu0 = -1.8105174530374e-09 wu0 = -8.95414305264101e-09 pu0 = 2.27821888296077e-15   a0 = 2.57551811198291 la0 = -9.26451720579159e-07 wa0 = -9.88634767548853e-06 pa0 = 5.48884995504779e-12   keta = 0.0805565649216189 lketa = -4.5849945136848e-08 wketa = -8.65031093894237e-07 pketa = 4.50623529463549e-13   a1 = 0.0   a2 = 1.54246581659637 la2 = -4.21244268350159e-07 wa2 = -3.66772476045626e-06 pa2 = 2.08785809718729e-12   ags = -2.45009036756156 lags = 1.78478452838403e-06 wags = 1.88517434172456e-05 pags = -1.01517066889696e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.147053561994433+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.1635084619579e-08 wvoff = -2.52666862140106e-07 pvoff = 2.67483830082796e-13   nfactor = {1.07112777586419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.87682393123814e-07 wnfactor = 4.80966456119758e-06 pnfactor = -3.15079829997579e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -54.6976859995376 letab = 3.07749182285744e-05 wetab = 0.000269156720183355 petab = -1.51437499312682e-10   dsub = 0.195324920036427 ldsub = 6.87261976223311e-08 wdsub = 1.41176517671706e-07 pdsub = -1.50019532385627e-13   voffl = 0.0   minv = 0.0   pclm = 1.64237004387538 lpclm = -5.74521059925369e-07 wpclm = -7.13657932101016e-06 ppclm = 4.02253468640667e-12   pdiblc1 = 0.644171048296386 lpdiblc1 = -3.13783392947467e-07 wpdiblc1 = 7.09465860942409e-07 ppdiblc1 = -5.84598682966564e-13   pdiblc2 = 0.00043   pdiblcb = 0.251698500472845 lpdiblcb = -2.6820869090904e-07 wpdiblcb = -6.50492050980012e-10 ppdiblcb = 3.65991546579808e-16   drout = -0.108059811559889 ldrout = 6.23436556256432e-07 wdrout = 3.48546326322919e-06 pdrout = -1.96105407949675e-12   pscbe1 = 800000000.0   pscbe2 = -4.83200297904129e-09 lpscbe2 = 1.91418529177648e-14 wpscbe2 = 9.36459327201553e-14 ppscbe2 = -1.30739178569451e-19   pvag = 0.0   delta = 0.01   alpha0 = 0.000328360992349073 lalpha0 = -1.84748315749498e-10 walpha0 = -1.61587780807945e-09 palpha0 = 9.09154258182204e-16   alpha1 = -6.3545624413236e-10 lalpha1 = 4.13795630286143e-16 walpha1 = 3.61921121362885e-15 palpha1 = -2.03630575881371e-21   beta0 = 162.608238578809 lbeta0 = -8.62116596830736e-05 wbeta0 = -0.000758930218585918 pbeta0 = 4.27094802434479e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 3215618293.13851 lbgidl = -1518.6895305036 wbgidl = -10199.8385011282 pbgidl = 0.00768525210892519   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.421220052079068 lkt1 = -4.90845098183373e-08 wkt1 = -6.90386254266983e-08 pkt1 = 3.88437541328274e-14   kt2 = -0.0367144850231195 lkt2 = -1.03939015195621e-08 wkt2 = -1.27222874502602e-08 pkt2 = 7.15804236643947e-15   at = 439285.019455141 lat = -0.199256938173075 wat = -2.28842420094424 pat = 1.24807916752632e-6   ute = -0.415425829980295 lute = -4.74285775017709e-08 wute = 1.29388998349895e-06 pute = -2.2381993658828e-13   ua1 = 3.2817400757718e-09 lua1 = -1.57660443518548e-15 wua1 = 1.30742661564253e-15 pua1 = -8.31421605017878e-22   ub1 = -2.72344529448287e-18 lub1 = 1.71734001132733e-24 wub1 = -2.01451368081573e-24 pub1 = 1.46102901889125e-30   uc1 = -5.34476908323868e-11 luc1 = 4.37550580345525e-17 wuc1 = 1.13321122309932e-17 puc1 = -6.37587696142163e-24   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.15 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.00214443219931+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.51434918816207e-09 wvth0 = -2.21685588604344e-07 pvth0 = 6.81200807407861e-14   k1 = 0.00103755770722369 lk1 = 2.58461915693318e-07 wk1 = 2.60642855712735e-07 pk1 = -8.83428253181225e-14   k2 = 0.168132919962517 lk2 = -8.96101507965653e-08 wk2 = -1.02488293498294e-07 pk2 = 4.14100763037387e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 70543.5223322177 lvsat = 0.00731073216162015 wvsat = 0.158522180185651 pvsat = -1.03902414153761e-7   ua = -3.94814505357321e-10 lua = -4.78276160266504e-16 wua = -5.76499364279383e-16 pua = 2.74615515812703e-23   ub = 1.08061958107146e-19 lub = 5.50910777464456e-25 wub = 2.03141131656479e-24 pub = -5.07758924494506e-31   uc = -3.62208260111838e-11 luc = 1.13367031901339e-17 wuc = 4.5736086243789e-17 puc = -1.41782921060887e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.010446337819473 lu0 = -1.63864599984193e-09 wu0 = -7.02563649643175e-09 pu0 = 1.19316781118827e-15   a0 = 1.31198782179594 la0 = -2.15541565168943e-07 wa0 = -5.78692231394371e-07 pa0 = 2.52009311293544e-13   keta = 0.0416161196304325 lketa = -2.39405708791055e-08 wketa = 2.62355715350357e-07 pketa = -1.83687130116212e-13   a1 = 0.0   a2 = 0.785980855071971 la2 = 4.38291743200976e-09 wa2 = 9.70270936548166e-08 pa2 = -3.0334356506053e-14   ags = -0.276422590269834 lags = 5.61796437504164e-07 wags = -2.74938990886524e-06 pags = 2.0019117633668e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.248903017975711+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.669289594815e-09 wvoff = 2.74221768418626e-07 pvoff = -2.89637352375084e-14   nfactor = {0.228229927566002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 8.61928752694611e-07 wnfactor = 4.16601698939911e-06 pnfactor = -2.78865771747425e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 2.39159688825581 leta0 = -1.06991067001448e-06 weta0 = -8.93454386494048e-06 peta0 = 5.02691389108238e-12   etab = 0.0171162692209475 letab = -9.70869031539364e-09 wetab = -7.58702171373926e-08 petab = 4.2986885069892e-14   dsub = 0.207451658361594 ldsub = 6.19032338245358e-08 wdsub = -3.78902158822502e-07 pdsub = 1.42596493999723e-13   voffl = 0.0   minv = 0.0   pclm = 0.183365767318676 lpclm = 2.46370188227942e-07 wpclm = 1.74945848462208e-06 ppclm = -9.77087852478647e-13   pdiblc1 = -0.500421881560025 lpdiblc1 = 3.30208083921085e-07 wpdiblc1 = 4.13488045068804e-07 ppdiblc1 = -4.18070316599067e-13   pdiblc2 = -0.0223768979208174 lpdiblc2 = 1.28320274323729e-08 wpdiblc2 = 7.42306350251015e-08 ppdiblc2 = -4.17649760292531e-14   pdiblcb = -0.25873232086764 lpdiblcb = 1.89790855483271e-08 wpdiblcb = -1.06480565856528e-06 ppdiblcb = 5.99100126123854e-13   drout = 2.523731747236 ldrout = -8.5730938280137e-07 wdrout = -5.9482993599131e-06 pdrout = 3.34673925526279e-12   pscbe1 = 800015319.568003 lpscbe1 = -0.00861937110175859 wpscbe1 = -0.0753882406243065 ppscbe1 = 4.24162889291202e-8   pscbe2 = 6.94922873163117e-08 lpscbe2 = -2.2675817125432e-14 wpscbe2 = -4.15368881061753e-13 ppscbe2 = 1.55651898227174e-19   pvag = 0.0   delta = 0.01   alpha0 = -8.80527474040498e-09 lalpha0 = 5.01044596939197e-15 walpha0 = -7.93724452551891e-15 palpha0 = 4.46579538534889e-21   alpha1 = 2.250552e-10 lalpha1 = -7.03608076176e-17   beta0 = 1.6822658135609 lbeta0 = 4.3314077816201e-06 wbeta0 = -1.12598175260384e-07 pbeta0 = 1.5517412186761e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = -168427457.348955 lbgidl = 385.303202459164 wbgidl = 3472.21377446176 pbgidl = -7.16403930819086e-6   cgidl = 509.73413487113 lcgidl = -0.000118004394175623 wcgidl = 0.000573839826670162 pcgidl = -3.22864092398047e-10   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.47338294432209 lkt1 = -1.97356844525086e-08 wkt1 = 1.93794629858882e-07 pkt1 = -1.09036222954542e-13   kt2 = 0.0395757132164887 lkt2 = -5.33176660766988e-08 wkt2 = -7.79437742069783e-08 pkt2 = 4.3854129232266e-14   at = -271.256318968022 lat = 0.0480541257159181 wat = 0.417094063447061 pat = -2.74148217714276e-7   ute = -0.476849762814122 lute = -1.28691387800119e-08 wute = 6.75031813998147e-07 pute = 1.24373186183312e-13   ua1 = 1.01453178257838e-09 lua1 = -3.00986895519715e-16 wua1 = -1.10008200473011e-15 pua1 = 5.23134230131348e-22   ub1 = 2.97352841063679e-19 lub1 = 1.77241899396863e-26 wub1 = 9.75786344256554e-25 pub1 = -2.21427406615377e-31   uc1 = -6.32076964459598e-11 luc1 = 4.92464080729619e-17 wuc1 = 4.8751062271753e-16 puc1 = -2.74292001744545e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.16 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.983076213462491+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.4710058128165e-10 wvth0 = -5.07839782237985e-08 pvth0 = 1.46897430746303e-14   k1 = 0.263452175081415 lk1 = 1.76421134546686e-07 wk1 = -8.5710372582091e-07 pk1 = 2.61107230439394e-13   k2 = 0.0874003555711931 lk2 = -6.43700833303906e-08 wk2 = 3.62090092388549e-07 pk2 = -1.03834781103152e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 127579.693995835 lvsat = -0.0105209424749498 wvsat = -0.792003169183225 pvsat = 1.93267930022226e-7   ua = -6.31916509581336e-10 lua = -4.04149063869918e-16 wua = -3.0756123509882e-15 pua = 8.08779237519938e-22   ub = -1.60383852362614e-19 lub = 6.34837138758101e-25 wub = 8.10861173123599e-24 pub = -2.40772270773648e-30   uc = 1.92401958179156e-13 luc = -4.74555757518327e-20 wuc = -2.07457751696567e-18 puc = 7.69138190746101e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00621132294166162 lu0 = -3.14619418472731e-10 wu0 = 3.67468111796053e-09 pu0 = -2.15215808714007e-15   a0 = 0.83420933474852 la0 = -6.61698545354108e-08 wa0 = 1.7345078983788e-06 pa0 = -4.7118495087848e-13   keta = -0.294979363468612 lketa = 8.12919677660135e-08 wketa = 6.93815261900249e-08 pketa = -1.23356065565504e-13   a1 = 0.0   a2 = 0.809136120402377 la2 = -2.85629841035832e-09 wa2 = 6.15597771144514e-07 pa2 = -1.92459255975075e-13   ags = 2.45826759610549 lags = -2.93171632983844e-07 wags = 1.63192571576998e-05 pags = -3.95967191822996e-12   b0 = 0.0   b1 = 1.79730994124424e-23 lb1 = -5.61907385410715e-30 wb1 = -1.24392579498309e-28 pb1 = 3.88898472691922e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.0919135995785685+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.0088293608412e-07 wvoff = -1.04434028675043e-06 pvoff = 3.83268868566434e-13   nfactor = {7.90025039991268+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.53663638373891e-06 wnfactor = -2.64675586681253e-05 pnfactor = 6.78856210894285e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -4.96587558741677 leta0 = 1.23031480983485e-06 weta0 = 3.03228511445592e-05 peta0 = -7.24643956989757e-12   etab = 0.148490346465222 letab = -5.07812190768893e-08 wetab = 1.89505744120486e-07 petab = -3.99797247058486e-14   dsub = 1.00117954454559 ldsub = -1.86246265056257e-07 wdsub = -8.41022944602491e-07 pdsub = 2.87073012224405e-13   voffl = 0.0   minv = 0.0   pclm = 2.14409314527263 lpclm = -3.66627697760824e-07 wpclm = -6.22373339604811e-06 ppclm = 1.51563491071032e-12   pdiblc1 = 1.87083628496936 lpdiblc1 = -4.11137326746331e-07 wpdiblc1 = -4.37078123242651e-06 ppdiblc1 = 1.07767406177851e-12   pdiblc2 = 0.0692896888584671 lpdiblc2 = -1.58264309251291e-08 wpdiblc2 = -2.67760625942309e-07 ppdiblc2 = 6.51544878170762e-14   pdiblcb = -0.624465996901287 lpdiblcb = 1.33321330556134e-07 wpdiblcb = 3.80287735201887e-06 ppdiblcb = -9.22722554939155e-13   drout = -4.59497231646062 ldrout = 1.36826801826461e-06 wdrout = 2.35092807259648e-05 pdrout = -5.8628196676259e-12   pscbe1 = 799945287.257133 lpscbe1 = 0.0132753905031677 wpscbe1 = 0.269243716524215 ppscbe1 = -6.53287568885136e-8   pscbe2 = -4.40683583949139e-08 lpscbe2 = 1.28275560284342e-14 wpscbe2 = 3.58809115974258e-13 ppscbe2 = -8.63855624101702e-20   pvag = 0.0   delta = 0.01   alpha0 = 3.19045526443035e-08 lalpha0 = -7.71699304450851e-15 walpha0 = 2.83473018768532e-14 palpha0 = -6.87813263279589e-21   alpha1 = -3.46625714285714e-10 lalpha1 = 1.08368370062857e-16   beta0 = 39.374359691844 lbeta0 = -7.45257306429856e-06 wbeta0 = 3.01676838899349e-06 pbeta0 = -8.23184782047654e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -5.60030200155297e-11 lagidl = 4.87724721716153e-17 wagidl = 7.67697444823869e-16 pagidl = -2.40011393754845e-22   bgidl = 2080244689.77566 lbgidl = -317.717160273581 wbgidl = 9907.30615088349 pbgidl = -0.00201901844968791   cgidl = -449.050481682606 lcgidl = 0.000181748110774504 wcgidl = -0.00204942795239344 pcgidl = 4.9726909951284e-10   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.53650925799 wkt1 = -1.54967270340524e-7   kt2 = -0.130965507226 wkt2 = 6.23274955435492e-8   at = 683537.132618207 lat = -0.165730361384622 wat = -2.95314318259109 pat = 7.79516014412599e-7   ute = -1.27370135609562 lute = 2.36256949640329e-07 wute = 4.79162546354378e-06 pute = -1.16263041922334e-12   ua1 = -2.35280509113946e-10 lua1 = 8.97519197303897e-17 wua1 = 2.56009703337911e-15 pua1 = -6.2117682398504e-22   ub1 = 2.20057783773615e-19 lub1 = 4.18895620607375e-26 wub1 = 1.19486406400433e-24 pub1 = -2.89919426761883e-31   uc1 = 9.43112490212e-11 wuc1 = -3.89836346443434e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.17 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.683057200844079+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -7.32431137649872e-08 wvth0 = -1.72957300413471e-06 pvth0 = 4.22027754743602e-13   k1 = -1.05598764433295 lk1 = 4.9656737344975e-07 wk1 = 1.32639271962858e-06 pk1 = -2.68691980091582e-13   k2 = 0.62979696421529 lk2 = -1.95976111658577e-07 wk2 = -4.13234397069731e-07 pk2 = 8.42884023700261e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 486833.779206231 lvsat = -0.0976896352022298 wvsat = -1.33419273368005 pvsat = 3.24823721572608e-7   ua = -1.088162183243e-09 lua = -2.93446526103997e-16 wua = 3.05561975042031e-15 pua = -6.78890657101618e-22   ub = 2.45081453021294e-18 lub = 1.26118560673381e-27 wub = -1.18089480120145e-23 pub = 2.42503415324635e-30   uc = -8.10393970488906e-13 luc = 1.95860822788329e-19 wuc = 7.86029704754329e-18 puc = -1.64143990383723e-24   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0103691835433468 lu0 = -1.32347439914443e-09 wu0 = -1.5818224732918e-08 pu0 = 2.57756160270536e-15   a0 = 1.39151042209027 la0 = -2.01392275765839e-07 wa0 = -1.95322595937297e-05 pa0 = 4.68894097987173e-12   keta = 0.375608276599924 lketa = -8.1418076044936e-08 wketa = -3.46149017055665e-06 pketa = 7.33367581189715e-13   a1 = 0.0   a2 = -3.57216130013436 la2 = 1.06021294511383e-06 wa2 = 1.88893287568163e-05 pa2 = -4.62636079487652e-12   ags = 1.25   b0 = 0.0   b1 = -4.19372319623654e-23 lb1 = 8.91744913001345e-30 wb1 = 2.9024935216272e-28 pb1 = -6.17180417451764e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.165721855004405+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.83707846550165e-08 wvoff = 5.18082190800868e-07 pvoff = 4.16580345834356e-15   nfactor = {-0.261706211471761+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 4.43764444534189e-07 wnfactor = 1.39242946395925e-05 pnfactor = -3.01203639393516e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -2.27049986671183 leta0 = 5.76314235714445e-07 weta0 = 8.80527859749781e-06 peta0 = -2.02545880222369e-12   etab = -0.314082520753951 letab = 6.14565362794365e-08 wetab = -1.70300808836236e-07 petab = 4.73230176904648e-14   dsub = 0.0464019091065495 ldsub = 4.54190708514017e-08 wdsub = 2.76696289973155e-06 pdsub = -5.88361457073117e-13   voffl = 0.0   minv = 0.0   pclm = 5.14987845450498 lpclm = -1.09594543362235e-06 wpclm = -1.60254131017913e-05 ppclm = 3.89389487115244e-12   pdiblc1 = 1.28840786884273 lpdiblc1 = -2.69818060714197e-07 wpdiblc1 = 5.71874744129926e-07 ppdiblc1 = -1.2160209906119e-13   pdiblc2 = 0.0480003877141518 lpdiblc2 = -1.06608374740747e-08 wpdiblc2 = -1.196765299343e-07 ppdiblc2 = 2.9223658929885e-14   pdiblcb = -1.83895350552948 lpdiblcb = 4.28002150674663e-07 wpdiblcb = 8.68048963954851e-06 ppdiblcb = -2.10621664516077e-12   drout = 1.35717084477475 ldrout = -7.59480940912125e-08 wdrout = -5.28582702797527e-06 pdrout = 1.12396768757461e-12   pscbe1 = 1145510168.95878 lpscbe1 = -83.8338963758215 wpscbe1 = -1700.27012197531 ppscbe1 = 0.000412550141855844   pscbe2 = 1.27029607036897e-08 lpscbe2 = -9.47323295012806e-16 wpscbe2 = -1.46660894741153e-14 ppscbe2 = 4.23371448941218e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 23.3531013287129 lbeta0 = -3.56520697758516e-06 wbeta0 = -4.18222843738638e-05 pbeta0 = 1.00564733022265e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.14782371605954e-09 lagidl = -2.43321639416168e-16 wagidl = -6.5240180636031e-15 pagidl = 1.52923587377886e-21   bgidl = -1978101156.34911 lbgidl = 666.991759138443 wbgidl = 18362.6114153157 pbgidl = -0.00407059680843924   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.499102860094567 lkt1 = -2.51278853107803e-07 wkt1 = -8.91255825751048e-07 pkt1 = 1.78651582507702e-13   kt2 = -0.19479594207674 lkt2 = 1.54876890513137e-08 wkt2 = 5.04100628789871e-07 pkt2 = -1.0719094950462e-13   at = -265284.086680194 lat = 0.0644897216235031 wat = 2.09904196250208 pat = -4.46336084822518e-7   ute = -0.3   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 4.93547947000197e-10 luc1 = -9.68699939242279e-17 wuc1 = -3.15297038094473e-15 puc1 = 6.70441315863325e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.18 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0785083674415+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.29965615015475e-8   k1 = 0.44156725201951 wk1 = -5.41497312046568e-8   k2 = 0.0186763023455965 wk2 = 5.60741270223443e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 316404.96230195 wvsat = -0.768137594089805   ua = -1.08000660920874e-09 wua = 2.60084264602229e-15   ub = 1.2344952447887e-18 wub = -2.45401319288716e-24   uc = -1.15543928775818e-11 wuc = -2.54287341855986e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.008619789691433 wu0 = 4.47027625295123e-9   a0 = 1.3692592466877 wa0 = -6.21031818558382e-7   keta = -0.0119692362598031 wketa = 3.49771639921365e-8   a1 = 0.0   a2 = 1.07010094796887 wa2 = -7.88976267277067e-7   ags = 0.249323491115106 wags = -3.00532481579464e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.226471217069939+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 4.37453441658362e-8   nfactor = {1.25272435765202+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.316004997689e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.341953277204447 wpclm = -5.64293730058397e-7   pdiblc1 = 0.39   pdiblc2 = 0.000134830687927477 wpdiblc2 = 1.66672658466809e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 862615051.653292 wpscbe1 = -308.13131154103   pscbe2 = 7.9142306921653e-09 wpscbe2 = 5.72235177942015e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.20031712910466e-10 walpha0 = -5.90681124570688e-16   alpha1 = 2.46052017904618e-10 walpha1 = -7.18728143503779e-16   beta0 = 1.48976041359756 wbeta0 = 2.39231717078135e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1819697250.51499 wbgidl = -1364.58458226916   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.423980008643474 wkt1 = -5.94148494127073e-8   kt2 = -0.0474262866831128 wkt2 = -1.53013868342091e-8   at = 90000.0   ute = -0.155175666687972 wute = -4.69292399763975e-8   ua1 = 1.73953927316707e-09 wua1 = 1.0817318179487e-15   ub1 = -7.7280610301252e-19 wub1 = 1.00285638556006e-25   uc1 = 1.1387738857419e-10 wuc1 = -9.57993346553485e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.19 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0785083674415+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.29965615015458e-8   k1 = 0.44156725201951 wk1 = -5.41497312046568e-8   k2 = 0.0186763023455965 wk2 = 5.60741270223446e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 316404.96230195 wvsat = -0.768137594089805   ua = -1.08000660920874e-09 wua = 2.60084264602229e-15   ub = 1.2344952447887e-18 wub = -2.45401319288716e-24   uc = -1.15543928775818e-11 wuc = -2.54287341855986e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00861978969143301 wu0 = 4.47027625295123e-9   a0 = 1.3692592466877 wa0 = -6.21031818558384e-7   keta = -0.0119692362598031 wketa = 3.49771639921365e-8   a1 = 0.0   a2 = 1.07010094796887 wa2 = -7.88976267277069e-7   ags = 0.249323491115106 wags = -3.00532481579464e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.226471217069939+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 4.37453441658366e-8   nfactor = {1.25272435765202+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.316004997689e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.341953277204447 wpclm = -5.64293730058398e-7   pdiblc1 = 0.39   pdiblc2 = 0.000134830687927477 wpdiblc2 = 1.66672658466809e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 862615051.653292 wpscbe1 = -308.13131154103   pscbe2 = 7.9142306921653e-09 wpscbe2 = 5.72235177942015e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.20031712910466e-10 walpha0 = -5.90681124570688e-16   alpha1 = 2.46052017904618e-10 walpha1 = -7.18728143503779e-16   beta0 = 1.48976041359756 wbeta0 = 2.39231717078135e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1819697250.51499 wbgidl = -1364.58458226916   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.423980008643474 wkt1 = -5.94148494127081e-8   kt2 = -0.0474262866831128 wkt2 = -1.53013868342091e-8   at = 90000.0   ute = -0.155175666687972 wute = -4.69292399763971e-8   ua1 = 1.73953927316707e-09 wua1 = 1.0817318179487e-15   ub1 = -7.7280610301252e-19 wub1 = 1.00285638556005e-25   uc1 = 1.1387738857419e-10 wuc1 = -9.57993346553504e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.20 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.07944380787821+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.54211761174215e-09 wvth0 = 5.83983952639036e-08 pvth0 = 3.70733498379238e-14   k1 = 0.528708250070802 lk1 = -7.02586322246271e-07 wk1 = -4.04856155152676e-07 pk1 = 2.82761894056741e-12   k2 = -0.0141519559745502 lk2 = 2.64682363005831e-07 wk2 = 1.42012419282648e-07 pk2 = -1.09978418944549e-12   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 540147.078990666 lvsat = -1.80395169221488 wvsat = -1.35163458227877 pvsat = 4.7045249898579e-6   ua = -1.60864139368819e-09 lua = 4.26219090146584e-15 wua = 4.42789085199611e-15 pua = -1.47308282933164e-20   ub = 1.69116573189314e-18 lub = -3.68196882280674e-24 wub = -4.2846109145625e-24 pub = 1.4759446753493e-29   uc = 3.20246884121063e-12 luc = -1.18979234054681e-16 wuc = -3.3706400641522e-16 puc = 6.67398281188534e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00697266921276628 lu0 = 1.32801361618765e-08 wu0 = 8.60103403814362e-09 pu0 = -3.3304804687688e-14   a0 = 1.36918459357151 la0 = 6.01901051403524e-10 wa0 = -5.31908129726297e-07 pa0 = -7.18572040277752e-13   keta = -0.0124041206201934 lketa = 3.50631516968859e-09 wketa = 6.5009582367067e-08 pketa = -2.42140517621613e-13   a1 = 0.0   a2 = 1.34443154173245 la2 = -2.21182826984086e-06 wa2 = -1.59030750841156e-06 pa2 = 6.46084371535812e-12   ags = 0.293502944889326 lags = -3.56202942819268e-07 wags = -9.41344359998847e-07 pags = 5.1666342017955e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.228966738385517+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.01204849887918e-08 wvoff = 6.11217260498661e-08 pvoff = -1.40099476880696e-13   nfactor = {1.16186927932755+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.32531606991886e-07 wnfactor = 1.72742371360156e-06 pnfactor = -3.31712017282785e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.201347706432053 lpclm = 1.13365181792119e-06 wpclm = -9.36646647530975e-07 ppclm = 3.00214678182527e-12   pdiblc1 = 0.39   pdiblc2 = 0.00032205401475534 lpdiblc2 = -1.50951390936875e-09 wpdiblc2 = -4.48776964278018e-10 ppdiblc2 = 4.96214751542811e-15   pdiblcb = -0.025   drout = 0.56   pscbe1 = 926210623.707949 lpscbe1 = -512.748075879614 wpscbe1 = -621.087805355135 ppscbe1 = 0.00252325491937238   pscbe2 = 6.40689415561773e-09 lpscbe2 = 1.21531088383568e-14 wpscbe2 = 1.11993444554345e-14 ppscbe2 = -4.41590092753547e-20   pvag = 0.0   delta = 0.01   alpha0 = 2.15202672236357e-10 lalpha0 = 3.89348068426177e-17 walpha0 = -5.6691721162788e-16 palpha0 = -1.91599827521371e-22   alpha1 = 2.47365326004197e-10 lalpha1 = -1.05887277893765e-17 walpha1 = -7.25190988083411e-16 palpha1 = 5.21075762958347e-23   beta0 = -9.21573971760501 lbeta0 = 8.63145721668389e-05 wbeta0 = 7.50116309440664e-05 pbeta0 = -4.11907752799663e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.53014491488423e-10 lagidl = -4.27436653625233e-16 wagidl = -2.60886549826069e-16 pagidl = 2.10343381031655e-21   bgidl = 1436107558.94081 lbgidl = 3092.74482369425 wbgidl = 801.808700833182 pbgidl = -0.0174668448072857   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.369649444339091 lkt1 = -4.38047672321961e-07 wkt1 = -1.92758458376714e-07 pkt1 = 1.07510124869034e-12   kt2 = -0.0433623137846803 lkt2 = -3.27663423218719e-08 wkt2 = -3.08423857355486e-08 pkt2 = 1.25301448299897e-13   at = 14407.7716211234 lat = 0.609472773032209 wat = 0.350392093041219 pat = -2.82508460425367e-6   ute = -0.0298010956067468 lute = -1.01084978103319e-06 wute = -4.59585131970809e-07 pute = 3.32709507571804e-12   ua1 = 1.2908175271376e-09 lua1 = 3.61788100096356e-15 wua1 = 2.18040301530058e-15 pua1 = -8.85818814527469e-21   ub1 = -6.20066700620844e-19 lub1 = -1.23148250982042e-24 wub1 = 2.0214170006898e-25 pub1 = -8.2122855208484e-31   uc1 = 3.61920815809313e-10 luc1 = -1.99988436207613e-15 wuc1 = -1.93098838991733e-17 puc1 = 7.84490681043677e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.21 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08515805003174+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.07570149258662e-08 wvth0 = 6.66706674674836e-08 pvth0 = 3.46610243730782e-15   k1 = 0.374270580034597 lk1 = -7.51619753257235e-08 wk1 = 6.31073200120606e-08 pk1 = 9.26452743751101e-13   k2 = 0.0449275604702652 lk2 = 2.46636744754988e-08 wk2 = -4.71910233598508e-08 pk2 = -3.31119093635257e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 96708.1393376625 lvsat = -0.00241980530087738 wvsat = -0.17968689021295 pvsat = -5.6674237940998e-8   ua = 1.60391840510412e-10 lua = -2.9247507390523e-15 wua = 2.39097293573291e-16 pua = 2.2867235912874e-21   ub = 1.44170029542897e-19 lub = 2.60291470339803e-24 wub = 2.847831124457e-25 pub = -3.8043470576035e-30   uc = -6.28245260991433e-11 luc = 1.49264544615809e-16 wuc = -1.2790793153154e-16 puc = -1.82327136564747e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0125602604811625 lu0 = -9.4202244535783e-09 wu0 = 2.39891478306094e-11 pu0 = 1.54062381140363e-15   a0 = 1.29744693422769 la0 = 2.9204604193268e-07 wa0 = -1.25981024894888e-07 pa0 = -2.36770692159583e-12   keta = -0.0137671797096042 lketa = 9.04393082257428e-09 wketa = 4.83526099539533e-08 pketa = -1.74469268531145e-13   a1 = 0.0   a2 = 0.8   ags = 0.110398086004728 lags = 3.87685814869937e-07 wags = -4.02980350595515e-08 pags = 1.50600916233678e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.217022426853907+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.84049289233664e-08 wvoff = -3.72131118493175e-08 pvoff = 2.59399372292371e-13   nfactor = {1.75211350170089+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.6654170001025e-06 wnfactor = -3.15640331534554e-08 pnfactor = 3.82901028867346e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.281737776899525 leta0 = -8.1958755846753e-07 weta0 = -5.89284559657696e-07 peta0 = 2.39404984487862e-12   etab = -0.246361959077213 letab = 7.1649479670153e-07 wetab = 5.15160724939212e-07 petab = -2.09291153724559e-12   dsub = 1.32127464809927 ldsub = -3.09278331380472e-06 wdsub = -2.22371537288812e-06 pdsub = 9.03415057507943e-12   voffl = 0.0   minv = 0.0   pclm = -0.01960736788749 lpclm = 2.03131229914459e-06 wpclm = 1.25360012223475e-06 ppclm = -5.89603297440222e-12   pdiblc1 = 0.39   pdiblc2 = -0.000867876264956714 lpdiblc2 = 3.32474206234007e-09 wpdiblc2 = 3.16312726731694e-09 ppdiblc2 = -9.71171186821039e-15   pdiblcb = 0.01064170425104 lpdiblcb = -1.44799342075037e-07 wpdiblcb = -1.75394330699287e-07 ppdiblcb = 7.12563672883491e-13   drout = 0.56   pscbe1 = 829306663.24877 lpscbe1 = -119.062363767655 wpscbe1 = -85.6060000908456 ppscbe1 = 0.000347786188997071   pscbe2 = 8.70478204734884e-09 lpscbe2 = 2.81762216967012e-15 wpscbe2 = 3.79556270326147e-15 ppscbe2 = -1.40801241852701e-20   pvag = 0.0   delta = 0.01   alpha0 = 2.78819688210145e-10 lalpha0 = -2.195180996991e-16 walpha0 = -8.79979231872964e-16 palpha0 = 1.08025783228308e-21   alpha1 = 3.94051622758831e-10 lalpha1 = -6.0652205106403e-16 walpha1 = -1.44704044457469e-15 palpha1 = 2.98472060851665e-21   beta0 = 13.3620740099792 lbeta0 = -5.41091183976648e-06 wbeta0 = -4.08624182538916e-05 pbeta0 = 5.88465626858302e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 8.27092575856233e-11 lagidl = -1.41811938772832e-16 wagidl = 8.50884730904776e-17 pagidl = 6.97862535164924e-22   bgidl = 2556208673.55055 lbgidl = -1457.82052836162 wbgidl = -4545.75120744717 pbgidl = 0.00425835528337059   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.504102658840388 lkt1 = 1.08187066133156e-07 wkt1 = 2.15219037771859e-07 pkt1 = -5.82363630307706e-13   kt2 = -0.0754354649697501 lkt2 = 9.75352604623377e-08 wkt2 = 8.45079739140203e-08 pkt2 = -3.43325306126108e-13   at = 173163.922121251 lat = -0.0354959967233305 wat = -0.312985006689432 pat = -1.30023590558137e-7   ute = -1.39520900355919 lute = 4.53630827131491e-06 wute = 6.30666993784774e-06 pute = -2.41617498886195e-11   ua1 = 3.61069113721713e-10 lua1 = 7.39511223574665e-15 wua1 = 1.24182606698556e-14 pua1 = -5.04508976912609e-20   ub1 = 4.43137385061683e-19 lub1 = -5.55089583006951e-24 wub1 = -8.62400725159857e-24 pub1 = 3.50362195726199e-29   uc1 = -5.39018932380831e-10 luc1 = 1.66030769463158e-15 wuc1 = 7.70670145951849e-16 puc1 = -3.13095382040953e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.22 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06773844154449+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.17333148504611e-09 wvth0 = 3.40193253756232e-09 pvth0 = 1.33966599315695e-13   k1 = 0.0959674454370201 lk1 = 4.98876645614353e-07 wk1 = 1.31939821968546e-06 pk1 = -1.66482060496945e-12   k2 = 0.151783658115618 lk2 = -1.95741773059515e-07 wk2 = -5.35183214500457e-07 pk2 = 6.7543214351462e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 235350.738043757 lvsat = -0.288389297810818 wvsat = -0.76199351511235 pvsat = 1.14441353422825e-6   ua = -1.73604329341946e-09 lua = 9.86908432726539e-16 wua = 4.42459154990813e-15 pua = -6.34643591061057e-21   ub = 1.66672490170332e-18 lub = -5.3756483300521e-25 wub = -3.31091624334954e-24 pub = 3.61227907023529e-30   uc = 5.20008470422209e-11 luc = -8.75786333897486e-17 wuc = -4.47142957842809e-16 puc = 4.76139159635875e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00586204269118676 lu0 = 4.39577409230175e-09 wu0 = 1.37983161119961e-08 pu0 = -2.68708264093089e-14   a0 = 2.79889840123788 la0 = -2.80490480907828e-06 wa0 = -5.68662880604956e-06 pa0 = 9.10189649642949e-12   keta = 0.104852257676451 lketa = -2.35625028268523e-07 wketa = -4.12986011644982e-07 pketa = 7.7710530324644e-13   a1 = 0.0   a2 = 0.8   ags = -1.42585992351966 lags = 3.5564299631193e-06 wags = 5.61635299304091e-06 pags = -1.01616142009623e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.280320106783758+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.0215527101178e-07 wvoff = 2.43571666927826e-07 pvoff = -3.19757982234959e-13   nfactor = {-0.665068359276642+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.32035415926046e-06 wnfactor = 7.15650569538841e-06 pnfactor = -1.09973754800667e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.759157133799049 leta0 = 1.32740183834595e-06 weta0 = 1.17856911931539e-06 peta0 = -1.25239233181107e-12   etab = -35.1331042133562 letab = 7.2675215066583e-05 wetab = 0.000172892950237616 petab = -3.57645890542094e-10   dsub = -0.643757896198541 ldsub = 9.60367483300625e-07 wdsub = 4.44743074577624e-06 pdsub = -4.72600891283017e-12   voffl = 0.0   minv = 0.0   pclm = 1.86392730800317 lpclm = -1.85373789766516e-06 wpclm = -4.88573767955113e-06 ppclm = 6.7671984703978e-12   pdiblc1 = 0.391279628332263 lpdiblc1 = -2.63941002400217e-09 wpdiblc1 = 3.94042961234308e-08 ppdiblc1 = -8.12767985474402e-14   pdiblc2 = 0.00107769315894229 lpdiblc2 = -6.88263363032114e-10 wpdiblc2 = -3.1873253678063e-09 ppdiblc2 = 3.38697305419495e-15   pdiblcb = -0.122061428134405 lpdiblcb = 1.28919181502214e-07 wpdiblcb = 3.50899199380092e-07 ppdiblcb = -3.7298936141238e-13   drout = 0.21088010504063 ldrout = 7.20107961899205e-07 wdrout = 4.00820616562778e-07 pdrout = -8.26747834905815e-13   pscbe1 = 741386673.50246 lpscbe1 = 62.2847480426926 wpscbe1 = 171.212000181689 ppscbe1 = -0.000181936377449071   pscbe2 = 1.33555134363087e-08 lpscbe2 = -6.77515312099122e-15 wpscbe2 = -7.45474782880296e-15 ppscbe2 = 9.1251938299662e-21   pvag = 0.0   delta = 0.01   alpha0 = 2.49322184351297e-10 lalpha0 = -1.58675427334693e-16 walpha0 = -7.3482077058891e-16 palpha0 = 7.80848474017059e-22   alpha1 = 1.0e-10   beta0 = 12.5772120818727 lbeta0 = -3.79202580210074e-06 wbeta0 = -2.50292429947905e-05 pbeta0 = 2.61884537357485e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -7.74764811249374e-11 lagidl = 1.88593252949641e-16 wagidl = 8.73369253123321e-16 pagidl = -9.28075356400459e-22   bgidl = 2580485906.4738 lbgidl = -1507.89567152398 wbgidl = -5232.57216191085 pbgidl = 0.00567501828324364   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.389986979026204 lkt1 = -1.27192271447411e-07 wkt1 = -3.24970257650686e-07 pkt1 = 5.31851337624059e-13   kt2 = -0.0112134329544985 lkt2 = -3.49315432095367e-08 wkt2 = -1.50053268525829e-07 pkt2 = 1.40489625857537e-13   at = 355783.540433254 lat = -0.412174160999163 wat = -1.07633880098295 pat = 1.44449895299585e-6   ute = 1.65439482048867 lute = -1.75392046111152e-06 wute = -9.87852305878628e-06 pute = 9.22244422357172e-12   ua1 = 3.55097550537859e-09 lua1 = 8.15490095872293e-16 wua1 = -1.22149136233953e-14 pua1 = 3.58423666621649e-22   ub1 = -6.06308777477555e-19 lub1 = -3.3862682962619e-24 wub1 = 3.88372570195038e-24 pub1 = 9.23729428877762e-30   uc1 = 7.24362546038596e-10 luc1 = -9.45590951252514e-16 wuc1 = -2.34822728453032e-15 puc1 = 3.30220253780534e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.23 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.12925378996215+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.01952153268022e-08 wvth0 = 2.22682286066155e-07 pvth0 = -9.90490369972268e-14   k1 = 0.609329347398712 lk1 = -4.66412191624156e-08 wk1 = -2.76581693203132e-07 pk1 = 3.11282977026633e-14   k2 = -0.0535912849815231 lk2 = 2.24974457233442e-08 wk2 = 1.21527548862592e-07 pk2 = -2.24136686439637e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -197081.568117857 lvsat = 0.171129703144147 wvsat = 0.829142151027175 pvsat = -5.46387687766924e-7   ua = 6.14894761022122e-11 lua = -9.23218194412433e-16 wua = -4.54795555014795e-15 pua = 3.18813359469882e-21   ub = 6.33558525271661e-19 lub = 5.6031701891338e-25 wub = 1.92009714532624e-24 pub = -1.94639453508037e-30   uc = -4.34590078900861e-11 luc = 1.38606359358083e-17 wuc = -3.63739087106242e-17 puc = 3.9640358804148e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0138851922596225 lu0 = -4.1299295188017e-09 wu0 = -2.43736389160425e-08 pu0 = 1.3692143537776e-14   a0 = -0.50781922538609 la0 = 7.0893899624216e-07 wa0 = 5.28688547853997e-06 pa0 = -2.55897677591816e-12   keta = -0.230120718341046 lketa = 1.20329985020758e-07 wketa = 6.6382492762269e-07 pketa = -3.67154919635081e-13   a1 = 0.0   a2 = 0.860689221267614 la2 = -6.44906727093749e-08 wa2 = -3.12673363871098e-07 pa2 = 3.32258598037255e-13   ags = 3.27596082210136 lags = -1.43990343036593e-06 wags = -9.3263961264458e-06 pags = 5.71711883787081e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.175804574906679+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -8.90690475101508e-09 wvoff = -1.11181914306198e-07 pvoff = 5.7216653820402e-14   nfactor = {3.2699697337517+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.61166849838981e-07 wnfactor = -6.01092950469745e-06 pnfactor = 2.99484152608217e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 70.6822077596497 letab = -3.9768156417788e-05 wetab = -0.000347843028037122 petab = 1.95707947939817e-10   dsub = 0.219652159591317 ldsub = 4.28751484362016e-08 wdsub = 2.14611452125829e-08 pdsub = -2.2805428426408e-14   voffl = 0.0   minv = 0.0   pclm = -0.449799147152498 lpclm = 6.04915755188546e-07 wpclm = 3.15907355757789e-06 ppclm = -1.78152365300251e-12   pdiblc1 = 1.08313617731787 lpdiblc1 = -7.37832469524968e-07 wpdiblc1 = -1.45070006330075e-06 ppdiblc1 = 1.50216471774235e-12   pdiblc2 = 0.000688708099695966 lpdiblc2 = -2.74913057644722e-10 wpdiblc2 = -1.27311347608566e-09 ppdiblc2 = 1.35285875800071e-15   pdiblcb = 0.251611239264651 lpdiblcb = -2.68159594437385e-07 wpdiblcb = -2.21075963034452e-10 ppdiblcb = 1.24385737689651e-16   drout = 0.76311834991874 ldrout = 1.3327861783842e-07 wdrout = -8.01641233125556e-07 pdrout = 4.51033820123296e-13   pscbe1 = 800000000.0   pscbe2 = 2.73877402911685e-08 lpscbe2 = -2.16863306015858e-14 wpscbe2 = -6.49087835857132e-14 ppscbe2 = 7.01780354786177e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.50742769378206 lbeta0 = 5.32681740491121e-07 wbeta0 = -5.93625166480933e-07 pbeta0 = 2.22237677909233e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.76772053628532e-10 lagidl = -1.87844701523716e-16 wagidl = -8.69902735686668e-16 pagidl = 9.2439170324461e-22   bgidl = 735750176.653581 lbgidl = 452.390614940724 wbgidl = 2003.69715052868 pbgidl = -0.00201451646638848   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.511056674771717 lkt1 = 1.46098790020919e-09 wkt1 = 3.73051185949302e-07 pkt1 = -2.09892773160144e-13   kt2 = -0.0315929944668784 lkt2 = -1.32754467231445e-08 wkt2 = -3.79253586044244e-08 pkt2 = 2.13382479144761e-14   at = -143039.19717653 lat = 0.117893835249023 wat = 0.577217843182151 pat = -3.12633172246464e-7   ute = 0.365626100165837 lute = -3.84425845685106e-07 wute = -2.54969952514162e-06 pute = 1.43455784142663e-12   ua1 = 8.85989090252241e-09 lua1 = -4.82596514391783e-15 wua1 = -2.61428890007621e-14 pua1 = 1.51588195656759e-20   ub1 = -8.61329217207105e-18 lub1 = 5.12225652420214e-24 wub1 = 2.69696713553339e-23 pub1 = -1.52947088284425e-29   uc1 = -3.79078280430305e-10 luc1 = 2.26967201704746e-16 wuc1 = 1.61377398525323e-15 puc1 = -9.07970567514908e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.24 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06131311266499+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.19692085336795e-08 wvth0 = 6.94859848855525e-08 pvth0 = -1.28549764935711e-14   k1 = 0.059244379978141 lk1 = 2.6285748673716e-07 wk1 = -2.57953730103472e-08 pk1 = -1.09973615917963e-13   k2 = 0.138406703036071 lk2 = -8.5527918258899e-08 wk2 = 4.37956744431017e-08 pk2 = 2.13212377156696e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 217657.063068969 lvsat = -0.0622180108295467 wvsat = -0.565429761971323 pvsat = 2.38251464218726e-7   ua = -7.90685635699103e-10 lua = -4.43752093858762e-16 wua = 1.37159917389423e-15 pua = -1.4243283612683e-22   ub = 9.23467378299504e-19 lub = 3.97203281663501e-25 wub = -1.98123316631053e-24 pub = 2.48642148798325e-31   uc = -5.44808491906469e-11 luc = 2.00619426814732e-17 wuc = 1.35594430882905e-16 puc = -5.71155638480763e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00898116841151265 lu0 = -1.37073934894886e-09 wu0 = 1.84523990290228e-10 pu0 = -1.25212123517246e-16   a0 = 0.54997619656988 la0 = 1.13783095623696e-07 wa0 = 3.17119913323367e-06 pa0 = -1.36861124196772e-12   keta = 0.133531166759215 lketa = -8.42743843082833e-08 wketa = -1.89962110385372e-07 pketa = 1.13218111855699e-13   a1 = 0.0   a2 = 0.678621557464772 la2 = 3.79475135173285e-08 wa2 = 6.25346727742194e-07 pa2 = -1.95507150267864e-13   ags = -3.69806964785218 lags = 2.48395112518779e-06 wags = 1.40886796550033e-05 pags = -7.45709256965217e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.199086820568669+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 4.1925713837559e-09 wvoff = 2.90741587350454e-08 pvoff = -2.16967426033774e-14   nfactor = {1.22535518972478+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.89210987983235e-07 wnfactor = -7.40878504370307e-07 pnfactor = 2.97105713601022e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.341633477020609 leta0 = 8.34766437560788e-08 weta0 = 1.15341259020392e-06 peta0 = -6.48953752927155e-13   etab = 0.0056199244666493 letab = -2.82239137631415e-09 wetab = -1.92962194557425e-08 petab = 9.09911738886661e-15   dsub = 0.286634281281112 ldsub = 5.18846145289871e-09 wdsub = -7.6856318771614e-07 pdsub = 4.21692282203942e-13   voffl = 0.0   minv = 0.0   pclm = 0.829425745391247 lpclm = -1.14824779902481e-07 wpclm = -1.42982993120411e-06 ppclm = 8.00367828118822e-13   pdiblc1 = -0.939030302559756 lpdiblc1 = 3.99915234380419e-07 wpdiblc1 = 2.57189859408384e-06 ppdiblc1 = -7.61102145651201e-13   pdiblc2 = -0.00568482040932858 lpdiblc2 = 3.31107627561583e-09 wpdiblc2 = -7.91178281460594e-09 ppdiblc2 = 5.08802639728708e-15   pdiblcb = -0.657309498062883 lpdiblcb = 2.43233751371105e-07 wpdiblcb = 8.96609450369387e-07 ppdiblcb = -5.04466547936932e-13   drout = 1.01871015778684 ldrout = -1.05270457568698e-08 wdrout = 1.45797539367733e-06 pdrout = -8.20312359547826e-13   pscbe1 = 800000000.0   pscbe2 = -5.04906866207438e-08 lpscbe2 = 2.21310317592788e-14 wpscbe2 = 1.75072396963997e-13 ppscbe2 = -6.48444959835103e-20   pvag = 0.0   delta = 0.01   alpha0 = -2.57802386628229e-08 lalpha0 = 1.45612057207734e-14 walpha0 = 7.55972692801772e-14 palpha0 = -4.25338963932604e-20   alpha1 = 4.0770095826472e-10 lalpha1 = -1.73124251756145e-16 walpha1 = -8.98807484071685e-16 palpha1 = 5.05703245223125e-22   beta0 = -10.4724583660738 lbeta0 = 1.12114868734363e-05 wbeta0 = 5.97013124420824e-05 pbeta0 = -3.37019854282977e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.24482110434344e-09 lagidl = -2.42041988331985e-15 wagidl = -2.03968395659247e-14 pagidl = 1.19109883875361e-20   bgidl = -138833525.395565 lbgidl = 944.464639894252 wbgidl = 3326.58078645522 pbgidl = -0.00275882106953891   cgidl = 666.047253142047 lcgidl = -0.000205952094413335 wcgidl = -0.000195383624754613 pcgidl = 1.09930251864686e-10   egidl = 2.41208050821963 legidl = -1.30086435298368e-06 wegidl = -1.13778457507463e-05 pegidl = 6.40160837750838e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.372249603050699 lkt1 = -7.66371453187609e-08 wkt1 = -3.03886810364636e-07 pkt1 = 1.70978267209938e-13   kt2 = 0.128659520116751 lkt2 = -1.03439601023449e-07 wkt2 = -5.1632894729982e-07 pkt2 = 2.90506286250876e-13   at = 67700.9690162429 lat = -0.000676590377346242 wat = 0.0825998741445795 pat = -3.43423073831024e-8   ute = -0.33967723176 lute = 1.24046103829828e-8   ua1 = 4.86802021878404e-10 lua1 = -1.1494716229004e-16 wua1 = 1.49689841787036e-15 pua1 = -3.92375147968623e-22   ub1 = 5.64932581426326e-19 lub1 = -4.17614946561167e-26 wub1 = -3.40984849933074e-25 pub1 = 7.13041575764605e-32   uc1 = 9.38881546460636e-12 luc1 = 8.40085180462481e-18 wuc1 = 1.30260124032831e-16 puc1 = -7.3289295665584e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.25 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.974819950539901+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.07184068678372e-09 wvth0 = -9.14133964801436e-08 pvth0 = 3.74482842978383e-14   k1 = 0.445195470783759 lk1 = 1.42194509609873e-07 wk1 = -1.75147015353924e-06 pk1 = 4.29537896117029e-13   k2 = 0.0393821196499728 lk2 = -5.4569070558236e-08 wk2 = 5.98389857726431e-07 pk2 = -1.52065978557664e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -129610.038868048 lvsat = 0.0463508813858384 wvsat = 0.473638359646669 pvsat = -8.66007151876802e-8   ua = -2.03246968439383e-09 lua = -5.55232124429389e-17 wua = 3.8165689256081e-15 pua = -9.06823289363152e-22   ub = 2.35748010453418e-18 lub = -5.11235890410563e-26 wub = -4.28190305451212e-24 pub = 9.67918981305894e-31   uc = 4.2679983996603e-11 luc = -1.03142258845222e-17 wuc = -2.11157761704011e-16 puc = 5.12923481379122e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00608840417901896 lu0 = -4.66351324830496e-10 wu0 = 4.27956953609658e-09 pu0 = -1.40547897286706e-15   a0 = 4.16249337981898 la0 = -1.01562705151294e-06 wa0 = -1.46441183409996e-05 pa0 = 4.20113398254164e-12   keta = -0.0673149705101581 lketa = -2.1482249644661e-08 wketa = -1.05096455899591e-06 pketa = 3.824001953844e-13   a1 = 0.0   a2 = 0.481649612352271 la2 = 9.95284284934109e-08 wa2 = 2.22717269718972e-06 pa2 = -6.96298817704e-13   ags = 14.6356646660369 lags = -3.24787090323786e-06 wags = -4.36062277095891e-05 pags = 1.05805278789993e-11   b0 = 0.0   b1 = -1.79730994124423e-23 lb1 = 5.61907385410714e-30 wb1 = 5.25001818485392e-29 pb1 = -1.64135518527636e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.103804859049946+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.55961905015348e-08 wvoff = -8.1201492520551e-08 pvoff = 1.27796164538699e-14   nfactor = {2.47292122532346+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.00825562254267e-07 wnfactor = 2.40557233319367e-07 pnfactor = -2.77123534799723e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.95369212969788 leta0 = -4.20514149299639e-07 weta0 = -3.7286335971197e-06 peta0 = 8.77359402985327e-13   etab = 0.0637725076777072 letab = -2.10030986862528e-08 wetab = 6.06405803886646e-07 petab = -1.86519111784851e-13   dsub = 0.14465787262736 ldsub = 4.95756819015904e-08 wdsub = 3.37395634812169e-06 pdsub = -8.73416740441323e-13   voffl = 0.0   minv = 0.0   pclm = -0.180918848434173 lpclm = 2.0104733322191e-07 wpclm = 5.21774874048917e-06 ppclm = -1.27791787264202e-12   pdiblc1 = 0.807505934928924 lpdiblc1 = -1.46118361835567e-07 wpdiblc1 = 8.61912292663274e-07 ppdiblc1 = -2.26495448347677e-13   pdiblc2 = 0.00631716031511607 lpdiblc2 = -4.41198974113099e-10 wpdiblc2 = 4.21298444602259e-08 ppdiblc2 = -1.05568878706618e-14   pdiblcb = 1.17773523857518 lpdiblcb = -3.30470965001948e-07 wpdiblcb = -5.06583098065298e-06 ppdiblcb = 1.35961890353704e-12   drout = 1.68921534252468 ldrout = -2.2015244570294e-07 wdrout = -7.4154719366211e-06 pdrout = 1.95386446690201e-12   pscbe1 = 800000000.0   pscbe2 = 5.87657914348052e-08 lpscbe2 = -1.2026695027052e-14 wpscbe2 = -1.47242074938913e-13 ppscbe2 = 3.59232558832718e-20   pvag = 0.0   delta = 0.01   alpha0 = 9.25294237957961e-08 lalpha0 = -2.24268905309644e-14 walpha0 = -2.69990247429205e-13 palpha0 = 6.55098936557273e-20   alpha1 = -9.98931993802571e-10 lalpha1 = 2.66642661112268e-16 walpha1 = 3.21002672882745e-15 palpha1 = -7.78874465429234e-22   beta0 = 83.6269549856618 lbeta0 = -1.82075655180236e-05 wbeta0 = -0.000214752120511406 pbeta0 = 5.21025869434149e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.49451318919219e-08 lagidl = 3.57908864152656e-15 wagidl = 7.40377289447136e-14 pagidl = -1.76128462424929e-20   bgidl = 8611617927.7977 lbgidl = -1791.25900152918 wbgidl = -22233.8571773736 pbgidl = 0.00523234313459661   cgidl = -1007.31161836445 lcgidl = 0.000317203476456714 wcgidl = 0.000697798659837903 pcgidl = -1.69312471225749e-10   egidl = -8.15743038649869 legidl = 2.00356639411927e-06 wegidl = 4.06351633955224e-05 pegidl = -9.85963477596276e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.940421003959704 lkt1 = 1.00994825118629e-07 wkt1 = 1.83269947665208e-06 pkt1 = -4.96999796390393e-13   kt2 = -0.51155276793557 lkt2 = 9.67150882886531e-08 wkt2 = 1.93521346627775e-06 pkt2 = -4.75939030845188e-13   at = 184488.770480255 lat = -0.037188895051452 wat = -0.497305132669341 pat = 1.46958034137188e-7   ute = -0.3   ua1 = 6.54531523711492e-11 lua1 = 1.67825055749691e-17 wua1 = 1.08017399425044e-15 pua1 = -2.62091257616937e-22   ub1 = 5.65342216226383e-19 lub1 = -4.18895620607373e-26 wub1 = -5.04295199098792e-25 pub1 = 1.22361178518933e-31   uc1 = 3.6259675067805e-11 wuc1 = -1.04162101242356e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.26 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.26685567284102+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.57871229009144e-08 wvth0 = 1.14332391285773e-06 pvth0 = -2.62145906965285e-13   k1 = -0.560403644911435 lk1 = 3.86191067843923e-07 wk1 = -1.11239705516949e-06 pk1 = 2.74474477674789e-13   k2 = 0.48684861236583 lk2 = -1.63141445417826e-07 wk2 = 2.9022047480191e-07 pk2 = -7.72923758236236e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -91439.4022728398 lvsat = 0.0370892344636504 wvsat = 1.51151399550671 pvsat = -3.38428783721488e-7   ua = -1.43461639592112e-10 lua = -5.13868346417538e-16 wua = -1.59329149124869e-15 pua = 4.05814422462155e-22   ub = -3.65505593942764e-19 lub = 6.09576214865993e-25 wub = 2.05028216766493e-24 pub = -5.6850977663271e-31   uc = 9.94738583000262e-13 luc = -1.9980130785648e-19 wuc = -1.02283642477066e-18 puc = 3.0563013800779e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00837972232482352 lu0 = -1.02231217709222e-09 wu0 = -6.02800212130122e-09 pu0 = 1.09552959894064e-15   a0 = -8.06858252800806 la0 = 1.9520967446104e-06 wa0 = 2.70212570296267e-05 pa0 = -5.9084693666364e-12   keta = -0.941351565245104 lketa = 1.90592241628637e-07 wketa = 3.01932478686806e-06 pketa = -6.05206670917342e-13   a1 = 0.0   a2 = 3.06557585704019 la2 = -5.27430267665177e-07 wa2 = -1.37752559061476e-05 pa2 = 3.18649845375257e-12   ags = 1.25   b0 = 0.0   b1 = 4.19372319623654e-23 lb1 = -8.91744913001346e-30 wb1 = -1.22500424313258e-28 pb1 = 2.60482452251226e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.189603193237908+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.7782542908359e-09 wvoff = 6.35603264040416e-07 pvoff = -1.6114445606857e-13   nfactor = {1.83591510232831+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.37363294170316e-08 wnfactor = 3.60181163476287e-06 pnfactor = -1.09269158025717e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.0900726594414918 leta0 = 3.16707517244315e-08 weta0 = -2.81119841986328e-06 peta0 = 6.54754766446184e-13   etab = -0.0762055740603547 letab = 1.2960903110507e-08 wetab = -1.34090330192258e-06 petab = 2.85972075030487e-13   dsub = 0.979643293338266 ldsub = -1.53023510608862e-07 wdsub = -1.82555733485914e-06 pdsub = 3.88182860569777e-13   voffl = 0.0   minv = 0.0   pclm = 1.79624423630145 lpclm = -2.78687563332171e-07 wpclm = 4.77962409352308e-07 ppclm = -1.27865596827637e-13   pdiblc1 = 1.52222643015005 lpdiblc1 = -3.19536713355029e-07 wpdiblc1 = -5.78756263206649e-07 ppdiblc1 = 1.23065488711489e-13   pdiblc2 = 0.0151528153037713 lpdiblc2 = -2.58506462925041e-09 wpdiblc2 = 4.19677600647381e-08 ppdiblc2 = -1.05175600371094e-14   pdiblcb = -0.182757519994824 lpdiblcb = -3.63723048038035e-10 wpdiblcb = 5.30279303261871e-07 ppdiblcb = 1.78989646850775e-15   drout = -0.764087114114552 ldrout = 3.75111955771091e-07 wdrout = 5.15297290480483e-06 pdrout = -1.09571785253189e-12   pscbe1 = 800000000.0   pscbe2 = 1.09272323885898e-08 lpscbe2 = -4.19242737196351e-16 wpscbe2 = -5.92765549977366e-15 ppscbe2 = 1.63500777939786e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 11.6121229994255 lbeta0 = -7.34030714547201e-07 wbeta0 = 1.59555654538452e-05 pbeta0 = -3.87586456382156e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.18858421541584e-09 lagidl = 2.41227426394477e-16 wagidl = 4.97354396360198e-15 pagidl = -8.552505270459e-22   bgidl = 2853624974.52647 lbgidl = -394.15110733336 wbgidl = -5414.51677356575 pbgidl = 0.00115133201769747   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.651665432951011 lkt1 = -2.85305843760514e-07 wkt1 = -1.64202268491821e-06 pkt1 = 3.46099839448698e-13   kt2 = -0.0491240579232608 lkt2 = -1.54876890513137e-08 wkt2 = -2.12756860482913e-07 pkt2 = 4.52401932993653e-14   at = -16838.4253221317 lat = 0.0116607330836475 wat = 0.876430378552149 pat = -1.86362402834572e-7   ute = -0.3   ua1 = 1.3462e-10   ub1 = 3.927e-19   uc1 = 2.40306869700692e-11 luc1 = 2.96721721405844e-18 wuc1 = -8.42456130708095e-16 puc1 = 1.79138186721508e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.27 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0569419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020595964   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.89624866e-10   ub = 3.9437962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01015016   a0 = 1.156653   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.14643813   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21149528+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7032502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.28 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0569419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020595964   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.89624866e-10   ub = 3.9437962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01015016   a0 = 1.156653   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.14643813   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21149528+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7032502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.29 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05945149305855+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.02339403584009e-8   k1 = 0.390108350640155 lk1 = 2.6543082607408e-7   k2 = 0.0344650819041385 lk2 = -1.11821677040387e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 77423.6776379675 lvsat = -0.193387835979627   ua = -9.27814543842969e-11 lua = -7.80813370542408e-16   ub = 2.2435675715032e-19 lub = 1.37083279488062e-24   uc = -1.1218922471776e-10 luc = 1.09500272742083e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.009917177867295 lu0 = 1.87845059646838e-9   a0 = 1.1870892682365 la0 = -2.45396612861797e-7   keta = 0.00985149156064635 lketa = -7.93889328420016e-08 wketa = -3.10192729707385e-25 pketa = 1.59251295241492e-29   a1 = 0.0   a2 = 0.8   ags = -0.028760239120425 lags = 1.41256102840836e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.208042108796165+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.78416693685451e-8   nfactor = {1.75324167155165+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.03063138208254e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.119307245944525 lpclm = 2.16141744959377e-06 ppclm = 8.07793566946316e-28   pdiblc1 = 0.39   pdiblc2 = 0.000168418108955 lpdiblc2 = 1.89245360671276e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 713585210.30066 lpscbe1 = 351.072008394549   pscbe2 = 1.02409176611441e-08 lpscbe2 = -2.96444381985355e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.1122212998938e-11 lalpha0 = -2.66581611471535e-17   alpha1 = -8.99142096746873e-13 lalpha1 = 7.2499656385495e-18 walpha1 = -3.37790056652293e-34 palpha1 = -1.61465456330906e-39   beta0 = 16.4640094294858 lbeta0 = -5.46993963405875e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.3701659983945e-11 lagidl = 2.92660375550365e-16   bgidl = 1710601607.95975 lbgidl = -2886.91709535839 wbgidl = -1.81898940354586e-12   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.435639062146295 lkt1 = -6.99936782063215e-8   kt2 = -0.0539210060677115 lkt2 = 1.01298021774776e-8   at = 134362.249869065 lat = -0.357676761559818   ute = -0.18713710806518 lute = 1.28159807982006e-7   ua1 = 2.0372644683357e-09 lua1 = 5.85337292668387e-16   ub1 = -5.508647904023e-19 lub1 = -1.51262481994686e-24   uc1 = 3.55310201317275e-10 luc1 = -1.97302782843743e-15 wuc1 = 1.97215226305253e-31   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.30 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.062333776056+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.1943612790595e-8   k1 = 0.39587496493943 lk1 = 2.42003159690503e-7   k2 = 0.0287720173015117 lk2 = -8.86928164493009e-08 wk2 = -1.32348898008484e-23 pk2 = -5.04870979341448e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 35193.488774603 lvsat = -0.0218218659561456   ua = 2.4224526035258e-10 lua = -2.14190563284761e-15   ub = 2.4166369548367e-19 lub = 1.30052096954389e-24   uc = -1.06612983359891e-10 luc = 8.68460227044348e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01256847301155 lu0 = -8.89280180579747e-9   a0 = 1.25431814105418 la0 = -5.18523186268071e-7   keta = 0.00278602515472579 lketa = -5.06845005335853e-8   a1 = 0.0   a2 = 0.8   ags = 0.09660231302358 lags = 9.03258360291149e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22976209622579+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.0398776922571e-8   nfactor = {1.7413077580682+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.54579967801672e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.40955456692973 lpclm = 1.2843351861936e-8   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -0.0494034161855245 lpdiblcb = 9.91422459251269e-8   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.00041685140221e-08 lpscbe2 = -2.00261773828812e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.2435539075844e-11 lalpha0 = 1.50301217626435e-16 palpha0 = -4.70197740328915e-38   alpha1 = -1.01333361605547e-10 lalpha1 = 4.15277842315342e-16 walpha1 = 7.70371977754894e-33 palpha1 = 5.28972457870029e-38   beta0 = -0.626911925893801 lbeta0 = 1.47348302127893e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1183874879615e-10 lagidl = 9.70968093325268e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.43042380621311 lkt1 = -9.11813751402025e-8   kt2 = -0.046504703916719 lkt2 = -1.99999487606265e-8   at = 66015.51916787 lat = -0.080008736237377   ute = 0.76383886567315 lute = -3.73531132001434e-6   ua1 = 4.6123807414194e-09 lua1 = -9.87642793277983e-15   ub1 = -2.50923600125864e-18 lub1 = 6.44352847938412e-24 wub1 = -1.46936793852786e-39   uc1 = -2.7518496724611e-10 luc1 = 5.88445802184582e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.31 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.066573811832+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.06892717035329e-8   k1 = 0.5476549354998 lk1 = -7.10639752261963e-8   k2 = -0.0314328714163614 lk2 = 3.54880748059554e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -25512.838357964 lvsat = 0.103393311227918   ua = -2.21312848954079e-10 lua = -1.18575306138354e-15   ub = 5.3325403183724e-19 lub = 6.99075661348239e-25   uc = -1.01075667170004e-10 luc = 7.54245439131587e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01058580741872 lu0 = -4.80328041273379e-9   a0 = 0.852117623456039 la0 = 3.11070884949521e-7   keta = -0.0365308458079778 lketa = 3.04119715551837e-8   a1 = 0.0   a2 = 0.8   ags = 0.49686238190986 lags = 7.766673232369e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.19693491401666+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.31181653490427e-9   nfactor = {1.78491531278+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.44526567237312e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.35568158 leta0 = 8.9865338280804e-07 peta0 = 2.01948391736579e-28   etab = 24.055684718764 letab = -4.9762554076942e-05 wetab = 4.97631856511901e-21 petab = 1.12081357413801e-26   dsub = 0.878791400000001 ldsub = -6.575512557132e-7   voffl = 0.0   minv = 0.0   pclm = 0.19132645357144 lpclm = 4.62968951143052e-7   pdiblc1 = 0.40476943553992 lpdiblc1 = -3.04639989831893e-8   pdiblc2 = -1.34671700000001e-05 lpdiblc2 = 4.7124506659446e-10   pdiblcb = -0.00193334529462572 lpdiblcb = 1.22867384286521e-9   drout = 0.34809846380408 ldrout = 4.37076160816079e-7   pscbe1 = 800000000.0   pscbe2 = 1.08034284890926e-08 lpscbe2 = -3.65120173474758e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.23897782188604e-12 lalpha0 = 1.08643022914693e-16   alpha1 = 1.0e-10   beta0 = 4.0086118080422 lbeta0 = 5.17342280927105e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.2151586247192e-10 lagidl = -1.29127373065436e-16   bgidl = 789148498.917399 lbgidl = 434.910318490012   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.50123845552 lkt1 = 5.48836114768618e-8   kt2 = -0.062583203828 lkt2 = 1.31641761393783e-8   at = -12694.121746 lat = 0.0823407600779259   ute = -1.7274539795 lute = 1.40332397156792e-06 wute = -1.6940658945086e-21   ua1 = -6.3072156952e-10 lua1 = 9.38194131651594e-16 wua1 = 3.94430452610506e-31   ub1 = 7.2325972446e-19 lub1 = -2.23940039320725e-25   uc1 = -7.9537953766e-11 luc1 = 1.84896837593995e-16 puc1 = 7.05296610493373e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.32 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.053019942308+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.6286414900289e-8   k1 = 0.514643384558759 lk1 = -3.59846467573118e-8   k2 = -0.011987110669152 lk2 = 1.48242704970624e-08 wk2 = -3.30872245021211e-24 pk2 = -3.15544362088405e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 86769.911681776 lvsat = -0.0159226057088111   ua = -1.4954738399868e-09 lua = 1.68218825805494e-16   ub = 1.2908914269758e-18 lub = -1.06018624947011e-25   uc = -5.59113814677852e-11 luc = 2.74312576831243e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00554103382327999 lu0 = 5.57487711177388e-10   a0 = 1.3021119966072 la0 = -1.67110235747081e-7   keta = -0.00286452614269639 lketa = -5.36313904129158e-9   a1 = 0.0   a2 = 0.753647507227639 la2 = 4.92559202146351e-8   ags = 0.0831291244128396 lags = 5.17315413603809e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21386698780376+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.0680848490072e-8   nfactor = {1.212166698692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.64097874539931e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -48.3996144876024 letab = 2.72312001611129e-5   dsub = 0.22699924455044 ldsub = 3.50678567694095e-8   voffl = 0.0   minv = 0.0   pclm = 0.63168935636104 lpclm = -4.97740315148235e-9   pdiblc1 = 0.586498346032599 lpdiblc1 = -2.2357604497131e-7   pdiblc2 = 0.000252865893758079 lpdiblc2 = 1.88229432388701e-10   pdiblcb = 0.25153555533135 lpdiblcb = -2.6811701178052e-07 wpdiblcb = -7.44462551297725e-23 ppdiblcb = 2.99767143983984e-29   drout = 0.48868163239184 ldrout = 2.8768714371432e-7   pscbe1 = 800000000.0   pscbe2 = 5.16663592447599e-09 lpscbe2 = 2.33866824253147e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.3042039380688 lbeta0 = 6.0876337940385e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.10335500312401e-11 lagidl = 1.28614849538097e-16   bgidl = 1421703002.1652 lbgidl = -237.266133732223   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.38334500188 lkt1 = -7.03944523122407e-8   kt2 = -0.044576496932 lkt2 = -5.97043486317338e-9   at = 54567.616988 lat = 0.0108658805531057   ute = -0.50724712472 lute = 1.06685799818211e-7   ua1 = -8.99589150400004e-11 lua1 = 3.63559186020276e-16   ub1 = 6.1960126416e-19 lub1 = -1.13788620384454e-25   uc1 = 1.7338685864e-10 luc1 = -8.38706792114924e-17 puc1 = 9.4039548065783e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.33 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.037525032888+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.75683900540385e-8   k1 = 0.0504135000235997 lk1 = 2.25208727017782e-7   k2 = 0.153399870352552 lk2 = -7.82287297310271e-08 wk2 = -2.64697796016969e-23 pk2 = -6.31088724176809e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24085.8226495999 lvsat = 0.0193458447760744   ua = -3.211274848808e-10 lua = -4.92513058738637e-16   ub = 2.452049532272e-19 lub = 4.82324321269954e-25   uc = -8.06096834027599e-12 luc = 5.08796941888806e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00904433901215999 lu0 = -1.41360491368368e-9   a0 = 1.63561581288 la0 = -3.54752155927177e-7   keta = 0.068498860692096 lketa = -4.55148922832455e-08 pketa = 1.89326617253043e-29   a1 = 0.0   a2 = 0.89270498554472 la2 = -2.898310127073e-8   ags = 1.125099170114 lags = -6.89365289694007e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.18913346942056+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.23516882601495e-9   nfactor = {0.971720201373598+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.9938221089816e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.736496854962879 leta0 = -1.38688497482605e-7   etab = -0.000986012091111663 letab = 2.92632908123304e-10   dsub = 0.02352161973992 ldsub = 1.49552100637551e-7   voffl = 0.0   minv = 0.0   pclm = 0.33993266952808 lpclm = 1.5917599561484e-7   pdiblc1 = -0.05855736927456 lpdiblc1 = 1.3935681257768e-7   pdiblc2 = -0.00839336834287296 lpdiblc2 = 5.05292937081832e-09 wpdiblc2 = 2.48154183765908e-24 ppdiblc2 = -3.94430452610506e-31   pdiblcb = -0.3503610224916 lpdiblcb = 7.05328749726289e-8   drout = 1.51783865160912 ldrout = -2.91355703264052e-7   pscbe1 = 800000000.0   pscbe2 = 9.44422187321678e-09 lpscbe2 = -6.80641604961539e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.96590176514319 lbeta0 = -3.26170962625641e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.73790566554872e-09 lagidl = 1.65723034286862e-15 wagidl = 7.88860905221012e-31 pagidl = -3.76158192263132e-37   bgidl = 1000000000.0   cgidl = 599.158926518552 lcgidl = -0.000168318180098545   egidl = -1.4830517670848 legidl = 8.90685080129057e-07 wegidl = 2.11758236813575e-22 pegidl = -5.04870979341448e-29   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.47628329704 lkt1 = -1.81038358000086e-8   kt2 = -0.048102372368 lkt2 = -3.98664335961322e-9   at = 95978.5043919999 lat = -0.0124334583141061   ute = -0.33967723176 lute = 1.2404610382983e-8   ua1 = 9.99255562559999e-10 lua1 = -2.49274269227633e-16 wua1 = -7.88860905221012e-31   ub1 = 4.48198612319999e-19 lub1 = -1.73509751585003e-26   uc1 = 5.39825306916e-11 luc1 = -1.66892669432604e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.34 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.00611473857143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.74833845949436e-9   k1 = -0.154409065411999 lk1 = 2.89244044230437e-7   k2 = 0.244237036749914 lk2 = -1.06627879759166e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 32537.0056514284 lvsat = 0.0167036838247486   ua = -7.25891872677145e-10 lua = -3.65968330066764e-16   ub = 8.91598148254288e-19 lub = 2.80237245563077e-25   uc = -2.96085169035249e-11 luc = 7.2453794296058e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00755348727028572 lu0 = -9.47508006807586e-10   a0 = -0.850826297999999 la0 = 4.22604132734124e-7   keta = -0.427105924230686 lketa = 1.09429996465443e-7   a1 = 0.0   a2 = 1.244107853178 la2 = -1.38844991001863e-7   ags = -0.292646780332859 lags = 3.74304729486404e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.131603667475429+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.12211710465369e-8   nfactor = {2.55527444614285+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.95697021078011e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.677218411817428 leta0 = -1.20155803574497e-7   etab = 0.271371632362262 letab = -8.48567163384906e-08 wetab = -2.91581165924942e-23 petab = 3.30335504061299e-29   dsub = 1.29971011669343 ldsub = -2.49432918673e-7   voffl = 0.0   minv = 0.0   pclm = 1.60534385618857 lpclm = -2.36439626960322e-7   pdiblc1 = 1.10257606183886 lpdiblc1 = -2.23657621058757e-7   pdiblc2 = 0.0207400414567257 lpdiblc2 = -4.05528160210861e-9   pdiblcb = -0.556519398572126 lpdiblcb = 1.34985817353692e-7   drout = -0.849423755746857 ldrout = 4.48740481246906e-7   pscbe1 = 800000000.0   pscbe2 = 8.35841459550001e-09 lpscbe2 = 2.71400455194675e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.1079484778457 lbeta0 = -3.70580162791528e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.04012081728377e-08 lagidl = -2.45055592933684e-15 pagidl = -3.00926553810506e-36   bgidl = 1000000000.0   cgidl = -768.424737566257 lcgidl = 0.000259240441473601 pcgidl = 5.16987882845642e-26   egidl = 5.75375631101714 legidl = -1.37181612379258e-6   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.313008131714287 lkt1 = -6.91498569371091e-8   kt2 = 0.150955108971428 lkt2 = -6.62195762106095e-8   at = 14239.5585142857 lat = 0.0131212422472108   ute = -0.3   ua1 = 4.35243768285714e-10 lua1 = -7.29427498893092e-17   ub1 = 3.927e-19   uc1 = 6.0045e-13   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.35 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.857830786089288+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.82309832028672e-08 wvth0 = -5.14550421942903e-08 pvth0 = 1.24849485279384e-14   k1 = 1.08647176599512 lk1 = -1.18407989405246e-08 wk1 = -5.92298962856989e-06 pk1 = 1.43714235749694e-12   k2 = -0.276305867352738 lk2 = 1.96756094064938e-08 wk2 = 2.51942691517889e-06 pk2 = -6.11308707845175e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1825500.85044608 lvsat = -0.418337477548537 wvsat = -4.08794937756393 pvsat = 9.91891861073358e-7   ua = -5.77355132519719e-09 lua = 8.58785664173797e-16 wua = 1.48524380701885e-14 pua = -3.60376586847439e-21   ub = 1.01682068559621e-17 lub = -1.97062053805772e-24 wub = -2.87191364211724e-23 pub = 6.96835382296043e-30   uc = -6.22082009881073e-13 luc = 2.12168839881864e-19 wuc = 3.69996475686474e-18 puc = -8.97752048676146e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00299889130580482 lu0 = 1.57610048822131e-10 wu0 = 9.68963235632139e-09 pu0 = -2.35107301567311e-15   a0 = -2.62595531921213 la0 = 8.53317888182993e-07 wa0 = 1.11231132738656e-05 pa0 = -2.6988899585442e-12   keta = -0.631480860028142 lketa = 1.59019122137466e-07 wketa = 2.11417938038556e-06 pketa = -5.12980256497991e-13   a1 = 0.0   a2 = -1.65029435741534 la2 = 5.63446972572081e-7   ags = -14.8979847726361 lags = 3.91811472926288e-06 wags = 4.71689449658275e-05 pags = -1.14449784686184e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.821289940828709+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.46122926947357e-07 wvoff = 2.4807869109339e-06 pvoff = -6.01933174495179e-13   nfactor = {3.33639467953319+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -3.85226472267372e-07 wnfactor = -7.81152530490725e-07 pnfactor = 1.89537287693209e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -1.54946890380923 leta0 = 4.20123153314524e-07 weta0 = 1.97797167504605e-06 peta0 = -4.79931091289823e-13   etab = -0.346097177894856 letab = 6.49646808446762e-08 wetab = -5.52538537696313e-07 petab = 1.34066845709558e-13   dsub = 0.358745919896382 ldsub = -2.11192478905583e-08 wdsub = -1.18899051662353e-08 pdsub = 2.88494280972537e-15   voffl = 0.0   minv = 0.0   pclm = 3.21738511047237 lpclm = -6.27582092817236e-07 wpclm = -3.67325005624586e-06 ppclm = 8.91270047147384e-13   pdiblc1 = 1.32409294779 lpdiblc1 = -2.7740603523217e-7   pdiblc2 = 0.0295202078956133 lpdiblc2 = -6.18568362650743e-9   pdiblcb = -0.340963036008864 lpdiblcb = 8.26836526540675e-08 wpdiblcb = 9.92404291811659e-07 ppdiblcb = -2.40794992556597e-13   drout = 1.0   pscbe1 = 546782850.815643 lpscbe1 = 61.4401026437945 wpscbe1 = 739.657978531206 ppscbe1 = -0.000179469132594856   pscbe2 = 5.35646802961673e-09 lpscbe2 = 9.99786766047454e-16 wpscbe2 = 1.03447822790425e-14 ppscbe2 = -2.51003728262232e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 17.934840186017 lbeta0 = -2.26968151307879e-06 wbeta0 = -2.51335826685395e-06 pbeta0 = 6.09836223152902e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.17273810446863e-09 lagidl = 3.57723247496219e-16 wagidl = 4.92725680481928e-15 pagidl = -1.19553973660774e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.111445859757879 lkt1 = -1.18056523480068e-07 wkt1 = 5.87057604381019e-07 pkt1 = -1.42442483011801e-13   kt2 = -0.0952722106735244 lkt2 = -6.47547182659724e-09 wkt2 = -7.79561588473442e-08 pkt2 = 1.89151264704017e-14   at = 118295.846023329 lat = -0.0121267672414085 wat = 0.481697469285807 pat = -1.1687811055257e-7   ute = 0.892372301693591 lute = -2.8931483053833e-07 wute = -3.48296981135811e-06 pute = 8.4510082908831e-13   ua1 = 1.40883460760295e-10 lua1 = -1.51975359195647e-18 wua1 = -1.82958331988667e-17 pua1 = 4.43926437570633e-24   ub1 = 2.69745542031596e-19 lub1 = 2.98334237725376e-26 wub1 = 3.59155160403834e-25 pub1 = -8.71446898100658e-32   uc1 = -6.93788001603463e-10 luc1 = 1.68485025120161e-16 wuc1 = 1.25432255056385e-15 puc1 = -3.04346315023711e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.36 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0569419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020595964   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.89624866e-10   ub = 3.9437962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01015016   a0 = 1.156653   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.14643813   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21149528+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7032502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.37 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0569419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020595964   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.89624866e-10   ub = 3.9437962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01015016   a0 = 1.156653   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.14643813   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21149528+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7032502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.38 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05945149305855+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.02339403584077e-8   k1 = 0.390108350640155 lk1 = 2.6543082607408e-7   k2 = 0.0344650819041385 lk2 = -1.11821677040387e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 77423.6776379675 lvsat = -0.193387835979627   ua = -9.27814543842973e-11 lua = -7.80813370542408e-16   ub = 2.24356757150319e-19 lub = 1.37083279488062e-24   uc = -1.12189224717759e-10 luc = 1.09500272742083e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.009917177867295 lu0 = 1.87845059646843e-9   a0 = 1.1870892682365 la0 = -2.4539661286179e-7   keta = 0.00985149156064634 lketa = -7.93889328420016e-08 wketa = 5.84196307615576e-24 pketa = -4.95503256091948e-29   a1 = 0.0   a2 = 0.8   ags = -0.0287602391204249 lags = 1.41256102840837e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.208042108796165+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.7841669368546e-8   nfactor = {1.75324167155165+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.0306313820826e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.119307245944525 lpclm = 2.16141744959377e-6   pdiblc1 = 0.39   pdiblc2 = 0.000168418108955 lpdiblc2 = 1.89245360671279e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 713585210.30066 lpscbe1 = 351.072008394549   pscbe2 = 1.02409176611441e-08 lpscbe2 = -2.9644438198535e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.1122212998938e-11 lalpha0 = -2.66581611471535e-17   alpha1 = -8.99142096746874e-13 lalpha1 = 7.2499656385495e-18 walpha1 = 8.89614124702307e-35 palpha1 = -5.71030245251134e-39   beta0 = 16.4640094294859 lbeta0 = -5.46993963405875e-05 pbeta0 = 1.03397576569128e-25   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37016599839449e-11 lagidl = 2.92660375550366e-16   bgidl = 1710601607.95975 lbgidl = -2886.91709535839   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.435639062146295 lkt1 = -6.99936782063198e-8   kt2 = -0.0539210060677116 lkt2 = 1.01298021774771e-8   at = 134362.249869065 lat = -0.357676761559819   ute = -0.18713710806518 lute = 1.28159807982005e-7   ua1 = 2.0372644683357e-09 lua1 = 5.85337292668381e-16   ub1 = -5.50864790402299e-19 lub1 = -1.51262481994686e-24   uc1 = 3.55310201317275e-10 luc1 = -1.97302782843743e-15 puc1 = 1.50463276905253e-36   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.39 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.062333776056+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.19436127905933e-8   k1 = 0.395874964939431 lk1 = 2.42003159690505e-7   k2 = 0.0287720173015117 lk2 = -8.86928164493009e-08 wk2 = -2.64697796016969e-23   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 35193.4887746031 lvsat = -0.0218218659561455   ua = 2.4224526035258e-10 lua = -2.1419056328476e-15 pua = 1.50463276905253e-36   ub = 2.4166369548367e-19 lub = 1.30052096954389e-24   uc = -1.06612983359891e-10 luc = 8.68460227044346e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01256847301155 lu0 = -8.89280180579744e-9   a0 = 1.25431814105418 la0 = -5.18523186268069e-7   keta = 0.00278602515472579 lketa = -5.06845005335853e-8   a1 = 0.0   a2 = 0.8   ags = 0.0966023130235798 lags = 9.03258360291148e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22976209622579+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.03987769225706e-8   nfactor = {1.7413077580682+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.54579967801672e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.40955456692973 lpclm = 1.28433518619368e-8   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -0.0494034161855245 lpdiblcb = 9.91422459251269e-8   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.00041685140221e-08 lpscbe2 = -2.00261773828812e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.24355390758441e-11 lalpha0 = 1.50301217626435e-16 palpha0 = -9.4039548065783e-38   alpha1 = -1.01333361605547e-10 lalpha1 = 4.15277842315342e-16 walpha1 = -2.77333911991762e-32 palpha1 = -1.93956567885677e-37   beta0 = -0.626911925893801 lbeta0 = 1.47348302127894e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1183874879615e-10 lagidl = 9.70968093325268e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.43042380621311 lkt1 = -9.11813751402042e-8   kt2 = -0.0465047039167189 lkt2 = -1.99999487606267e-8   at = 66015.5191678701 lat = -0.0800087362373769   ute = 0.76383886567315 lute = -3.73531132001433e-06 wute = -4.2351647362715e-22 pute = -8.07793566946316e-28   ua1 = 4.6123807414194e-09 lua1 = -9.87642793277982e-15   ub1 = -2.50923600125864e-18 lub1 = 6.44352847938411e-24   uc1 = -2.7518496724611e-10 luc1 = 5.88445802184582e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.40 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.066573811832+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.06892717035337e-8   k1 = 0.5476549354998 lk1 = -7.10639752261963e-8   k2 = -0.0314328714163614 lk2 = 3.54880748059554e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -25512.838357964 lvsat = 0.103393311227918   ua = -2.21312848954079e-10 lua = -1.18575306138353e-15   ub = 5.33254031837239e-19 lub = 6.9907566134824e-25   uc = -1.01075667170004e-10 luc = 7.54245439131587e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01058580741872 lu0 = -4.80328041273379e-9   a0 = 0.85211762345604 la0 = 3.11070884949519e-7   keta = -0.0365308458079778 lketa = 3.04119715551837e-8   a1 = 0.0   a2 = 0.8   ags = 0.49686238190986 lags = 7.76667323236895e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.196934914016659+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.31181653490427e-9   nfactor = {1.78491531278+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.44526567237314e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.35568158 leta0 = 8.9865338280804e-07 weta0 = 2.11758236813575e-22 peta0 = -2.01948391736579e-28   etab = 24.055684718764 letab = -4.97625540769419e-05 wetab = 5.29395592033938e-21 petab = -2.70610844927016e-26   dsub = 0.878791400000001 ldsub = -6.575512557132e-07 wdsub = -1.6940658945086e-21   voffl = 0.0   minv = 0.0   pclm = 0.191326453571439 lpclm = 4.62968951143052e-7   pdiblc1 = 0.404769435539919 lpdiblc1 = -3.04639989831901e-8   pdiblc2 = -1.34671700000003e-05 lpdiblc2 = 4.7124506659446e-10   pdiblcb = -0.00193334529462572 lpdiblcb = 1.22867384286521e-09 wpdiblcb = -3.30872245021211e-24   drout = 0.34809846380408 ldrout = 4.3707616081608e-7   pscbe1 = 800000000.0   pscbe2 = 1.08034284890926e-08 lpscbe2 = -3.65120173474757e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.2389778218861e-12 lalpha0 = 1.08643022914693e-16   alpha1 = 1.0e-10   beta0 = 4.00861180804218 lbeta0 = 5.17342280927106e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.2151586247192e-10 lagidl = -1.29127373065436e-16   bgidl = 789148498.917398 lbgidl = 434.91031849001   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.501238455519999 lkt1 = 5.48836114768618e-8   kt2 = -0.062583203828 lkt2 = 1.31641761393783e-8   at = -12694.1217460001 lat = 0.082340760077926   ute = -1.7274539795 lute = 1.40332397156792e-6   ua1 = -6.3072156952e-10 lua1 = 9.38194131651594e-16   ub1 = 7.2325972446e-19 lub1 = -2.23940039320725e-25   uc1 = -7.95379537660001e-11 luc1 = 1.84896837593995e-16 wuc1 = 4.93038065763132e-32 puc1 = 1.41059322098675e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.41 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.053019942308+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.62864149002886e-8   k1 = 0.514643384558759 lk1 = -3.59846467573116e-8   k2 = -0.011987110669152 lk2 = 1.48242704970624e-08 wk2 = -6.61744490042422e-24 pk2 = 1.26217744835362e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 86769.9116817759 lvsat = -0.0159226057088111   ua = -1.4954738399868e-09 lua = 1.68218825805494e-16   ub = 1.2908914269758e-18 lub = -1.06018624947011e-25   uc = -5.59113814677852e-11 luc = 2.74312576831244e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00554103382327999 lu0 = 5.57487711177388e-10   a0 = 1.3021119966072 la0 = -1.67110235747082e-7   keta = -0.00286452614269639 lketa = -5.36313904129159e-9   a1 = 0.0   a2 = 0.753647507227639 la2 = 4.92559202146355e-8   ags = 0.0831291244128396 lags = 5.17315413603808e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21386698780376+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.06808484900718e-8   nfactor = {1.212166698692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.64097874539931e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -48.3996144876024 letab = 2.72312001611128e-5   dsub = 0.22699924455044 ldsub = 3.50678567694095e-8   voffl = 0.0   minv = 0.0   pclm = 0.63168935636104 lpclm = -4.97740315148277e-9   pdiblc1 = 0.5864983460326 lpdiblc1 = -2.2357604497131e-7   pdiblc2 = 0.000252865893758079 lpdiblc2 = 1.88229432388702e-10   pdiblcb = 0.251535555331349 lpdiblcb = -2.6811701178052e-07 wpdiblcb = 1.45583787809333e-22 ppdiblcb = 1.92482060873927e-28   drout = 0.48868163239184 ldrout = 2.8768714371432e-7   pscbe1 = 800000000.0   pscbe2 = 5.16663592447599e-09 lpscbe2 = 2.33866824253147e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.3042039380688 lbeta0 = 6.08763379403857e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.10335500312401e-11 lagidl = 1.28614849538097e-16   bgidl = 1421703002.1652 lbgidl = -237.266133732224   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.38334500188 lkt1 = -7.03944523122405e-8   kt2 = -0.0445764969319999 lkt2 = -5.97043486317335e-9   at = 54567.616988 lat = 0.0108658805531057   ute = -0.507247124719999 lute = 1.06685799818211e-7   ua1 = -8.99589150400002e-11 lua1 = 3.63559186020275e-16   ub1 = 6.19601264159999e-19 lub1 = -1.13788620384454e-25   uc1 = 1.7338685864e-10 luc1 = -8.38706792114923e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.42 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.037525032888+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.75683900540385e-8   k1 = 0.0504135000236001 lk1 = 2.25208727017782e-7   k2 = 0.153399870352552 lk2 = -7.82287297310271e-08 wk2 = 1.05879118406788e-22 pk2 = 2.52435489670724e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24085.8226496 lvsat = 0.0193458447760744   ua = -3.21127484880799e-10 lua = -4.92513058738635e-16   ub = 2.452049532272e-19 lub = 4.82324321269955e-25   uc = -8.06096834027601e-12 luc = 5.08796941888812e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00904433901216001 lu0 = -1.41360491368368e-9   a0 = 1.63561581288 la0 = -3.54752155927178e-7   keta = 0.068498860692096 lketa = -4.55148922832455e-08 wketa = 5.29395592033938e-23 pketa = -2.52435489670724e-29   a1 = 0.0   a2 = 0.89270498554472 la2 = -2.898310127073e-8   ags = 1.125099170114 lags = -6.89365289694002e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.18913346942056+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.23516882601501e-9   nfactor = {0.971720201373596+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.99382210898159e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.73649685496288 leta0 = -1.38688497482605e-7   etab = -0.000986012091111663 letab = 2.92632908123304e-10   dsub = 0.02352161973992 ldsub = 1.49552100637551e-7   voffl = 0.0   minv = 0.0   pclm = 0.33993266952808 lpclm = 1.5917599561484e-7   pdiblc1 = -0.0585573692745607 lpdiblc1 = 1.3935681257768e-7   pdiblc2 = -0.00839336834287296 lpdiblc2 = 5.05292937081832e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = -2.36658271566304e-30   pdiblcb = -0.3503610224916 lpdiblcb = 7.05328749726288e-8   drout = 1.51783865160912 ldrout = -2.91355703264052e-7   pscbe1 = 800000000.0   pscbe2 = 9.44422187321677e-09 lpscbe2 = -6.8064160496157e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.96590176514319 lbeta0 = -3.26170962625638e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.73790566554872e-09 lagidl = 1.65723034286862e-15 wagidl = -1.57772181044202e-30 pagidl = -1.31655367292096e-36   bgidl = 1000000000.0   cgidl = 599.158926518552 lcgidl = -0.000168318180098545 wcgidl = -8.67361737988404e-19   egidl = -1.4830517670848 legidl = 8.90685080129058e-07 wegidl = 4.2351647362715e-22 pegidl = -1.0097419586829e-28   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.47628329704 lkt1 = -1.81038358000081e-8   kt2 = -0.0481023723680001 lkt2 = -3.98664335961318e-9   at = 95978.5043919999 lat = -0.0124334583141061   ute = -0.33967723176 lute = 1.24046103829831e-8   ua1 = 9.99255562559999e-10 lua1 = -2.49274269227633e-16   ub1 = 4.4819861232e-19 lub1 = -1.73509751584999e-26   uc1 = 5.39825306916e-11 luc1 = -1.66892669432604e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.43 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.00611473857143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.74833845949394e-9   k1 = -0.154409065412001 lk1 = 2.89244044230437e-7   k2 = 0.244237036749914 lk2 = -1.06627879759166e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 32537.0056514284 lvsat = 0.0167036838247487   ua = -7.25891872677145e-10 lua = -3.65968330066761e-16   ub = 8.91598148254291e-19 lub = 2.80237245563078e-25   uc = -2.96085169035249e-11 luc = 7.2453794296058e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00755348727028572 lu0 = -9.47508006807586e-10   a0 = -0.850826297999998 la0 = 4.22604132734123e-7   keta = -0.427105924230685 lketa = 1.09429996465443e-07 wketa = 4.2351647362715e-22   a1 = 0.0   a2 = 1.244107853178 la2 = -1.38844991001863e-7   ags = -0.292646780332859 lags = 3.74304729486403e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.131603667475429+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.1221171046537e-8   nfactor = {2.55527444614285+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.95697021078011e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.677218411817428 leta0 = -1.20155803574497e-7   etab = 0.271371632362262 letab = -8.48567163384905e-08 wetab = 2.60561892954204e-23 petab = 4.4866463984445e-29   dsub = 1.29971011669343 ldsub = -2.49432918673e-7   voffl = 0.0   minv = 0.0   pclm = 1.60534385618857 lpclm = -2.36439626960322e-7   pdiblc1 = 1.10257606183886 lpdiblc1 = -2.23657621058757e-7   pdiblc2 = 0.0207400414567257 lpdiblc2 = -4.05528160210861e-9   pdiblcb = -0.556519398572126 lpdiblcb = 1.34985817353692e-7   drout = -0.849423755746855 ldrout = 4.48740481246906e-7   pscbe1 = 800000000.0   pscbe2 = 8.35841459550002e-09 lpscbe2 = 2.71400455194675e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.1079484778457 lbeta0 = -3.70580162791524e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.04012081728377e-08 lagidl = -2.45055592933684e-15   bgidl = 1000000000.0   cgidl = -768.424737566257 lcgidl = 0.000259240441473602 wcgidl = -4.33680868994202e-19 pcgidl = -1.03397576569128e-25   egidl = 5.75375631101714 legidl = -1.37181612379258e-6   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.313008131714286 lkt1 = -6.91498569371093e-8   kt2 = 0.150955108971428 lkt2 = -6.62195762106096e-8   at = 14239.5585142856 lat = 0.0131212422472107   ute = -0.3   ua1 = 4.35243768285714e-10 lua1 = -7.29427498893091e-17   ub1 = 3.927e-19   uc1 = 6.0045e-13   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.44 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.25338225871071+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.77448350110456e-08 wvth0 = 7.08416028983582e-07 pvth0 = -1.7188864844052e-13   k1 = -6.97133921903205 lk1 = 1.9432903428445e-06 wk1 = 9.55640531329095e-06 pk1 = -2.31874707240629e-12   k2 = 3.28426725519255 lk2 = -8.4425473190165e-07 wk2 = -4.32058430941638e-06 pk2 = 1.04833793566817e-12   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3907730.48029061 lvsat = 0.972762306078754 wvsat = 6.92582995114342 pvsat = -1.68046952768554e-6   ua = 1.52692659846084e-08 lua = -4.24700144224281e-15 wua = -2.55717019888386e-14 pua = 6.20466662716782e-21   ub = -3.42061235057744e-17 lub = 8.79627823225329e-24 wub = 5.65258248004647e-23 pub = -1.37153130779351e-29   uc = 8.64823990997546e-13 luc = -1.48611058359322e-19 wuc = 8.43555581743671e-19 puc = -2.04678639243121e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0011056135222581 lu0 = 6.16991183666335e-10 wu0 = 1.33266988748371e-08 pu0 = -3.23356356159273e-15   a0 = 11.6312274140987 la0 = -2.60601641586208e-06 wa0 = -1.62655364099359e-05 pa0 = 3.94663722343402e-12   keta = 2.83623676817464 lketa = -6.82380947734399e-07 wketa = -4.54745252107589e-06 pketa = 1.10338478480881e-12   a1 = 0.0   a2 = -1.65029435741533 la2 = 5.63446972572082e-7   ags = 51.7124524144875 lags = -1.22441085289464e-05 wags = -8.07925158310864e-05 pags = 1.96033344562231e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {3.91680826482956+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.00351974547716e-06 wvoff = -6.62129968987993e-06 pvoff = 1.60657891415309e-12   nfactor = {6.89059980608302+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.24761169576316e-06 wnfactor = -7.60893056604925e-06 pnfactor = 1.84621569468506e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.188921131794713 leta0 = -1.67632814434523e-09 weta0 = -1.36154894340863e-06 peta0 = 3.30363512530782e-13   etab = -1.88691963219585 letab = 4.38826759511361e-07 wetab = 2.40744641972347e-06 petab = -5.84137984388863e-13   dsub = 0.341955385747058 ldsub = -1.70452262656341e-08 wdsub = 2.03654194951626e-08 pdsub = -4.94142465546735e-15   voffl = 0.0   minv = 0.0   pclm = -0.671947704916299 lpclm = 3.16117842843042e-07 wpclm = 3.79832241196061e-06 ppclm = -9.21617353393298e-13   pdiblc1 = 1.32409294779 lpdiblc1 = -2.7740603523217e-7   pdiblc2 = 0.0295202078956134 lpdiblc2 = -6.18568362650743e-9   pdiblcb = 1.06134355415248 lpdiblcb = -2.57569213769501e-07 wpdiblcb = -1.70148584522639e-06 ppdiblcb = 4.12845122514041e-13   drout = 1.0   pscbe1 = 1591303591.20113 lpscbe1 = -192.000320761856 wpscbe1 = -1266.91044252454 ppscbe1 = 0.000307400615953269   pscbe2 = 1.15967643403723e-08 lpscbe2 = -5.1434625020164e-16 wpscbe2 = -1.64309027442319e-15 ppscbe2 = 3.98676138005475e-22   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 19.8953099678517 lbeta0 = -2.74536598000359e-06 wbeta0 = -6.27950344958301e-06 pbeta0 = 1.52364615799993e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.15871250886701e-09 lagidl = -1.42116526642231e-15 wagidl = -9.15676921061436e-15 pagidl = 2.22178016772505e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.194147429333331 lkt1 = -1.92205067958581e-7   kt2 = -0.135852349333335 lkt2 = 3.3708118575416e-9   at = 841975.085197033 lat = -0.187718850476037 wat = -0.908520888430771 pat = 2.20441691327066e-7   ute = -0.920690322000002 lute = 1.50603058349436e-7   ua1 = 1.18283012314007e-09 lua1 = -2.54335607858461e-16 wua1 = -2.01991934177957e-15 pua1 = 4.90109189250712e-22   ub1 = -6.67261694100266e-20 lub1 = 1.11474246893311e-25 wub1 = 1.00553151718943e-24 pub1 = -2.43980156267808e-31   uc1 = -4.08494297366666e-11 luc1 = 1.00573159195453e-17 wuc1 = 1.23259516440783e-32 puc1 = -2.93873587705572e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.45 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0569419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020595964   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.89624866e-10   ub = 3.9437962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01015016   a0 = 1.156653   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.14643813   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21149528+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7032502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.46 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0569419+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.42302944   k2 = 0.020595964   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 53438.0   ua = -1.89624866e-10   ub = 3.9437962e-19   uc = -9.8608028e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01015016   a0 = 1.156653   keta = 4.9707517e-6   a1 = 0.0   a2 = 0.8   ags = 0.14643813   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21149528+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7032502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.14877095   pdiblc1 = 0.39   pdiblc2 = 0.00019189   pdiblcb = -0.025   drout = 0.56   pscbe1 = 757128280.0   pscbe2 = 9.873241e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.7815831e-11   alpha1 = 6.3056523e-17   beta0 = 9.6797043   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 1352540500.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.4443203   kt2 = -0.052664618   at = 90000.0   ute = -0.17124159   ua1 = 2.1098632e-9   ub1 = -7.3847396e-19   uc1 = 1.1059776e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.47 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05945149305855+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.02339403583942e-8   k1 = 0.390108350640155 lk1 = 2.65430826074087e-7   k2 = 0.0344650819041386 lk2 = -1.11821677040387e-07 wk2 = 4.2351647362715e-22   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 77423.6776379663 lvsat = -0.193387835979625   ua = -9.27814543842957e-11 lua = -7.80813370542416e-16   ub = 2.24356757150324e-19 lub = 1.3708327948806e-24   uc = -1.1218922471776e-10 luc = 1.09500272742083e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00991717786729507 lu0 = 1.87845059646822e-9   a0 = 1.18708926823649 la0 = -2.45396612861756e-7   keta = 0.00985149156064633 lketa = -7.93889328420018e-08 wketa = 4.85968609874904e-23 pketa = -6.98141901120595e-29   a1 = 0.0   a2 = 0.8   ags = -0.0287602391204249 lags = 1.41256102840839e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.208042108796167+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.78416693685511e-8   nfactor = {1.75324167155165+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.0306313820826e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.11930724594453 lpclm = 2.16141744959378e-06 ppclm = -1.29246970711411e-26   pdiblc1 = 0.39   pdiblc2 = 0.000168418108954998 lpdiblc2 = 1.89245360671279e-10   pdiblcb = -0.025   drout = 0.56   pscbe1 = 713585210.300659 lpscbe1 = 351.07200839452   pscbe2 = 1.0240917661144e-08 lpscbe2 = -2.96444381985371e-15   pvag = 0.0   delta = 0.01   alpha0 = 2.11222129989381e-11 lalpha0 = -2.66581611471519e-17   alpha1 = -8.99142096746871e-13 lalpha1 = 7.2499656385495e-18 walpha1 = 4.60267164053168e-33 palpha1 = -3.92826334815807e-38   beta0 = 16.4640094294857 lbeta0 = -5.4699396340588e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37016599839457e-11 lagidl = 2.92660375550359e-16   bgidl = 1710601607.95975 lbgidl = -2886.91709535848   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.435639062146301 lkt1 = -6.99936782063164e-8   kt2 = -0.0539210060677116 lkt2 = 1.01298021774784e-8   at = 134362.249869063 lat = -0.357676761559816   ute = -0.18713710806518 lute = 1.28159807982002e-7   ua1 = 2.0372644683357e-09 lua1 = 5.85337292668305e-16   ub1 = -5.50864790402291e-19 lub1 = -1.51262481994687e-24   uc1 = 3.55310201317275e-10 luc1 = -1.97302782843744e-15 wuc1 = 3.15544362088405e-30   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.48 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.06233377605599+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.19436127906069e-8   k1 = 0.395874964939431 lk1 = 2.42003159690502e-7   k2 = 0.0287720173015115 lk2 = -8.86928164493013e-08 pk2 = -4.03896783473158e-28   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 35193.4887746028 lvsat = -0.021821865956146   ua = 2.42245260352582e-10 lua = -2.14190563284761e-15 pua = -1.20370621524202e-35   ub = 2.41663695483673e-19 lub = 1.3005209695439e-24   uc = -1.0661298335989e-10 luc = 8.68460227044354e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0125684730115501 lu0 = -8.89280180579776e-9   a0 = 1.25431814105418 la0 = -5.18523186268042e-7   keta = 0.00278602515472581 lketa = -5.06845005335849e-08 pketa = -4.03896783473158e-28   a1 = 0.0   a2 = 0.8   ags = 0.0966023130235811 lags = 9.03258360291143e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.229762096225791+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.03987769225714e-8   nfactor = {1.74130775806819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.54579967801639e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.409554566929728 lpclm = 1.28433518619368e-8   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -0.0494034161855241 lpdiblcb = 9.91422459251263e-8   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.00041685140221e-08 lpscbe2 = -2.00261773828853e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.2435539075844e-11 lalpha0 = 1.50301217626435e-16 palpha0 = 7.52316384526264e-37   alpha1 = -1.01333361605547e-10 lalpha1 = 4.15277842315343e-16 walpha1 = -7.39557098644699e-32 palpha1 = 1.36357344695385e-36   beta0 = -0.626911925893751 lbeta0 = 1.47348302127894e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1183874879615e-10 lagidl = 9.70968093325272e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.430423806213106 lkt1 = -9.11813751402042e-8   kt2 = -0.0465047039167201 lkt2 = -1.99999487606272e-8   at = 66015.5191678703 lat = -0.080008736237378   ute = 0.763838865673144 lute = -3.73531132001433e-06 wute = 3.3881317890172e-21 pute = 1.93870456067116e-26   ua1 = 4.61238074141942e-09 lua1 = -9.87642793277988e-15   ub1 = -2.50923600125864e-18 lub1 = 6.44352847938412e-24   uc1 = -2.7518496724611e-10 luc1 = 5.88445802184579e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.49 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.066573811832+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.06892717035219e-8   k1 = 0.547654935499807 lk1 = -7.1063975226192e-8   k2 = -0.0314328714163614 lk2 = 3.54880748059555e-08 pk2 = 4.03896783473158e-28   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -25512.8383579645 lvsat = 0.10339331122792   ua = -2.21312848954077e-10 lua = -1.18575306138355e-15   ub = 5.33254031837247e-19 lub = 6.9907566134823e-25   uc = -1.01075667170004e-10 luc = 7.54245439131602e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.01058580741872 lu0 = -4.80328041273393e-9   a0 = 0.852117623456039 la0 = 3.11070884949512e-7   keta = -0.0365308458079783 lketa = 3.04119715551836e-8   a1 = 0.0   a2 = 0.8   ags = 0.496862381909864 lags = 7.76667323236946e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.196934914016666+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.31181653490173e-9   nfactor = {1.78491531278002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.44526567237321e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.355681580000002 leta0 = 8.98653382808038e-07 weta0 = 1.6940658945086e-21 peta0 = 3.23117426778526e-27   etab = 24.0556847187639 letab = -4.97625540769422e-05 wetab = 1.55854062294791e-19 petab = -3.0049920690403e-25   dsub = 0.878791400000004 ldsub = -6.57551255713187e-7   voffl = 0.0   minv = 0.0   pclm = 0.191326453571435 lpclm = 4.62968951143066e-7   pdiblc1 = 0.404769435539926 lpdiblc1 = -3.04639989831884e-8   pdiblc2 = -1.34671700000033e-05 lpdiblc2 = 4.71245066594462e-10   pdiblcb = -0.00193334529462572 lpdiblcb = 1.2286738428652e-9   drout = 0.348098463804078 ldrout = 4.37076160816094e-7   pscbe1 = 800000000.0   pscbe2 = 1.08034284890924e-08 lpscbe2 = -3.65120173474777e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.23897782188558e-12 lalpha0 = 1.08643022914695e-16   alpha1 = 1.0e-10   beta0 = 4.00861180804225 lbeta0 = 5.17342280927124e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.21515862471924e-10 lagidl = -1.29127373065434e-16   bgidl = 789148498.917404 lbgidl = 434.910318490016   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.501238455520003 lkt1 = 5.48836114768576e-8   kt2 = -0.0625832038280008 lkt2 = 1.31641761393782e-8   at = -12694.1217460004 lat = 0.0823407600779258   ute = -1.72745397950001 lute = 1.40332397156792e-6   ua1 = -6.30721569519997e-10 lua1 = 9.38194131651599e-16 pua1 = 6.01853107621011e-36   ub1 = 7.23259724460002e-19 lub1 = -2.23940039320724e-25   uc1 = -7.95379537659998e-11 luc1 = 1.84896837593995e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.50 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05301994230801+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.62864149003038e-8   k1 = 0.514643384558767 lk1 = -3.59846467573065e-8   k2 = -0.011987110669152 lk2 = 1.48242704970622e-08 wk2 = -5.29395592033938e-23 pk2 = -7.57306469012171e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 86769.9116817759 lvsat = -0.0159226057088109   ua = -1.49547383998679e-09 lua = 1.68218825805489e-16   ub = 1.29089142697577e-18 lub = -1.06018624947011e-25   uc = -5.59113814677849e-11 luc = 2.74312576831245e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00554103382327997 lu0 = 5.57487711177375e-10   a0 = 1.30211199660721 la0 = -1.67110235747072e-7   keta = -0.0028645261426965 lketa = -5.36313904129147e-9   a1 = 0.0   a2 = 0.75364750722764 la2 = 4.92559202146389e-8   ags = 0.0831291244128494 lags = 5.17315413603813e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.213866987803762+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.06808484900727e-8   nfactor = {1.21216669869202+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.64097874539928e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -48.3996144876019 letab = 2.72312001611127e-5   dsub = 0.226999244550441 ldsub = 3.50678567694102e-8   voffl = 0.0   minv = 0.0   pclm = 0.631689356361036 lpclm = -4.97740315147854e-9   pdiblc1 = 0.586498346032599 lpdiblc1 = -2.2357604497131e-7   pdiblc2 = 0.000252865893758079 lpdiblc2 = 1.88229432388699e-10   pdiblcb = 0.251535555331349 lpdiblcb = -2.68117011780518e-07 wpdiblcb = -6.88214269644119e-22 ppdiblcb = -4.54383881407303e-28   drout = 0.488681632391845 ldrout = 2.87687143714317e-7   pscbe1 = 800000000.0   pscbe2 = 5.16663592447596e-09 lpscbe2 = 2.33866824253147e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.30420393806878 lbeta0 = 6.08763379403884e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.10335500312399e-11 lagidl = 1.28614849538095e-16   bgidl = 1421703002.16521 lbgidl = -237.266133732221   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.383345001879995 lkt1 = -7.03944523122417e-8   kt2 = -0.0445764969320006 lkt2 = -5.97043486317372e-9   at = 54567.6169880005 lat = 0.0108658805531059   ute = -0.507247124720003 lute = 1.06685799818208e-7   ua1 = -8.9958915040001e-11 lua1 = 3.63559186020272e-16   ub1 = 6.19601264160012e-19 lub1 = -1.13788620384454e-25   uc1 = 1.7338685864e-10 luc1 = -8.38706792114919e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.51 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.03752503288801+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.75683900540343e-8   k1 = 0.0504135000235948 lk1 = 2.25208727017785e-7   k2 = 0.153399870352552 lk2 = -7.82287297310267e-08 wk2 = -4.2351647362715e-22 pk2 = -1.0097419586829e-28   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24085.8226496 lvsat = 0.0193458447760744   ua = -3.21127484880785e-10 lua = -4.92513058738635e-16   ub = 2.45204953227184e-19 lub = 4.82324321269951e-25   uc = -8.06096834027601e-12 luc = 5.087969418888e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00904433901215995 lu0 = -1.41360491368365e-9   a0 = 1.63561581287999 la0 = -3.54752155927172e-7   keta = 0.0684988606920964 lketa = -4.55148922832454e-08 pketa = -1.0097419586829e-28   a1 = 0.0   a2 = 0.892704985544711 la2 = -2.89831012707334e-8   ags = 1.12509917011398 lags = -6.89365289694062e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.189133469420561+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.23516882601543e-9   nfactor = {0.971720201373586+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.99382210898156e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.736496854962873 leta0 = -1.38688497482606e-7   etab = -0.000986012091111661 letab = 2.92632908123306e-10   dsub = 0.0235216197399168 ldsub = 1.49552100637551e-7   voffl = 0.0   minv = 0.0   pclm = 0.339932669528082 lpclm = 1.5917599561484e-7   pdiblc1 = -0.0585573692745633 lpdiblc1 = 1.39356812577679e-7   pdiblc2 = -0.00839336834287298 lpdiblc2 = 5.05292937081832e-09 wpdiblc2 = -1.32348898008484e-23 ppdiblc2 = -6.31088724176809e-30   pdiblcb = -0.350361022491597 lpdiblcb = 7.05328749726285e-8   drout = 1.51783865160913 ldrout = -2.91355703264052e-7   pscbe1 = 800000000.0   pscbe2 = 9.44422187321693e-09 lpscbe2 = -6.80641604961255e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.96590176514314 lbeta0 = -3.26170962625604e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.73790566554872e-09 lagidl = 1.65723034286862e-15 wagidl = 1.89326617253043e-29 pagidl = -6.01853107621011e-36   bgidl = 1000000000.0   cgidl = 599.158926518554 lcgidl = -0.000168318180098544   egidl = -1.4830517670848 legidl = 8.90685080129053e-07 wegidl = 1.01643953670516e-20 pegidl = -2.42338070083895e-27   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.476283297039998 lkt1 = -1.81038358000103e-8   kt2 = -0.0481023723679996 lkt2 = -3.98664335961315e-9   at = 95978.5043919999 lat = -0.0124334583141059   ute = -0.33967723176 lute = 1.24046103829831e-8   ua1 = 9.99255562559982e-10 lua1 = -2.49274269227631e-16   ub1 = 4.48198612320005e-19 lub1 = -1.73509751584977e-26   uc1 = 5.39825306916001e-11 luc1 = -1.66892669432602e-17 wuc1 = -7.88860905221012e-31   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.52 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.00611473857137+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.74833845949309e-9   k1 = -0.154409065412011 lk1 = 2.89244044230432e-7   k2 = 0.244237036749919 lk2 = -1.06627879759165e-7   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 32537.0056514256 lvsat = 0.0167036838247494   ua = -7.25891872677086e-10 lua = -3.65968330066783e-16   ub = 8.91598148254198e-19 lub = 2.80237245563088e-25   uc = -2.96085169035249e-11 luc = 7.2453794296058e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0075534872702856 lu0 = -9.47508006807529e-10   a0 = -0.850826298000015 la0 = 4.22604132734121e-7   keta = -0.427105924230684 lketa = 1.09429996465444e-7   a1 = 0.0   a2 = 1.24410785317798 la2 = -1.38844991001863e-7   ags = -0.292646780332888 lags = 3.74304729486396e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.131603667475424+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.12211710465383e-8   nfactor = {2.55527444614279+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.95697021078016e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.677218411817421 leta0 = -1.20155803574498e-7   etab = 0.271371632362262 letab = -8.48567163384907e-08 wetab = 1.43267682094184e-21 petab = -1.51461293802434e-28   dsub = 1.29971011669342 ldsub = -2.49432918673001e-7   voffl = 0.0   minv = 0.0   pclm = 1.60534385618854 lpclm = -2.3643962696032e-7   pdiblc1 = 1.10257606183886 lpdiblc1 = -2.23657621058758e-7   pdiblc2 = 0.0207400414567256 lpdiblc2 = -4.05528160210864e-9   pdiblcb = -0.556519398572121 lpdiblcb = 1.34985817353692e-7   drout = -0.849423755746869 ldrout = 4.48740481246903e-7   pscbe1 = 800000000.0   pscbe2 = 8.35841459549965e-09 lpscbe2 = 2.71400455194662e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 10.1079484778456 lbeta0 = -3.70580162791585e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.04012081728378e-08 lagidl = -2.45055592933685e-15   bgidl = 1000000000.0   cgidl = -768.424737566254 lcgidl = 0.000259240441473599   egidl = 5.75375631101713 legidl = -1.37181612379257e-6   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.31300813171427 lkt1 = -6.91498569371102e-8   kt2 = 0.150955108971431 lkt2 = -6.62195762106094e-8   at = 14239.5585142821 lat = 0.0131212422472107   ute = -0.3   ua1 = 4.35243768285715e-10 lua1 = -7.29427498893089e-17   ub1 = 3.927e-19   uc1 = 6.0045e-13   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.53 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.25267182576442+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.75350911593783e-06 wvth0 = -1.13090933157435e-05 pvth0 = 2.74401578394536e-12   k1 = -1.00247386789329 lk1 = 4.95016791774881e-7   k2 = -3.11204936494495 lk2 = 7.07734740175272e-07 wk2 = 5.92018852398513e-06 pk2 = -1.4364627030827e-12   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7098581.44977881 lvsat = -1.69778720800942 wvsat = -10.6957399152612 pvsat = 2.59519294155913e-6   ua = -5.7596196205274e-09 lua = 8.55405303216141e-16 wua = 8.09643128395651e-15 pua = -1.96450189387666e-21   ub = 4.52096053080999e-17 lub = -1.04729953756875e-23 wub = -7.0622108374304e-23 pub = 1.71356071317244e-29   uc = 1.39170303375087e-12 luc = -2.76451935534899e-19   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.146421302368221 lu0 = -3.46421169265404e-08 wu0 = -2.19329851289619e-07 pu0 = 5.32177564572104e-14   a0 = 1.47188469974935 la0 = -1.40973818337785e-7   keta = -0.00407095205653363 lketa = 6.78563688705152e-9   a1 = 0.0   a2 = -1.65029435741531 la2 = 5.63446972572074e-7   ags = 1.25   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {16.6228040302068+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.08647714599673e-06 wvoff = -2.69641351032701e-05 pvoff = 6.54252381318722e-12   nfactor = {-59.2367327175559+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.47973920131075e-05 wnfactor = 9.82637193777294e-05 pnfactor = -2.38425123423734e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.661493019318002 leta0 = 2.04666460653341e-7   etab = -0.383245075882805 letab = 7.39781725166745e-8   dsub = 0.354675487375331 ldsub = -2.01316062845181e-8   voffl = 0.0   minv = 0.0   pclm = 1.70045847648271 lpclm = -2.5951804819924e-7   pdiblc1 = 1.32409294779001 lpdiblc1 = -2.77406035232168e-7   pdiblc2 = 0.0295202078956136 lpdiblc2 = -6.18568362650738e-9   pdiblcb = -0.00139285918277766 lpdiblcb = 2.91024089339606e-10   drout = 1.0   pscbe1 = 800000000.0   pscbe2 = 1.05705014008804e-08 lpscbe2 = -2.65335863089229e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 15.973175092467 lbeta0 = -1.79370701811001e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.39457132204014e-10 lagidl = -3.34565803395543e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.194147429333327 lkt1 = -1.92205067958573e-7   kt2 = -0.135852349333334 lkt2 = 3.37081185754117e-9   at = 274519.156533334 lat = -0.0500324788569344   ute = -0.920690321999984 lute = 1.50603058349433e-7   ua1 = -7.8797672666664e-11 lua1 = 5.1783237260494e-17   ub1 = 5.61321934000003e-19 lub1 = -4.09140888218893e-26   uc1 = -4.08494297366666e-11 luc1 = 1.00573159195453e-17 wuc1 = -4.93038065763132e-32 puc1 = -1.17549435082229e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.54 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.22018585571533+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.5646314332372e-7   k1 = 0.214861425044933 wk1 = 3.2704073618464e-7   k2 = 0.0520850050141133 wk2 = -4.94706122707028e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 47987.59018134 wvsat = 0.00856282383240919   ua = 3.44169001577158e-09 wua = -5.70494892075117e-15   ub = -1.64199871850573e-18 wub = 3.19923630495839e-24   uc = -2.7937238741136e-10 wuc = 2.83988436891214e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0260855438916973 wu0 = -2.50351605670567e-8   a0 = 0.783374013593332 wa0 = 5.864370400181e-7   keta = -0.0200886954067375 wketa = 3.15679974876172e-8   a1 = 0.0   a2 = 0.8   ags = -0.0656680853125332 wags = 3.33227815138276e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.319878220519267+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.70274173315858e-7   nfactor = {2.43585188798533+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.15094816761619e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.594026026461021 wpclm = -6.99514514884491e-7   pdiblc1 = 0.39   pdiblc2 = -0.000946599370666533 wpdiblc2 = 1.78861484556857e-9   pdiblcb = 0.580662666666666 wpdiblcb = -9.51521608297866e-7   drout = 0.56   pscbe1 = 627343825.1902 wpscbe1 = 203.896855410188   pscbe2 = 7.15160495793333e-09 wpscbe2 = 4.27580507512772e-15   pvag = 0.0   delta = 0.01   alpha0 = 7.17677495617133e-11 walpha0 = -8.47607408314149e-17   alpha1 = 2.5401143235454e-16 walpha1 = -2.99998220893157e-22   beta0 = -51.856518105586 wbeta0 = 9.66760022277611e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -4.14462774745333e-11 wagidl = 2.22218070945401e-16   bgidl = 2420143596.69 wbgidl = -1677.24951775067   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.137583350960667 wkt1 = -4.81896691240042e-7   kt2 = -0.05321158589764 wkt2 = 8.59309649237735e-10   at = 332265.066666667 wat = -0.380608643319147   ute = 3.12434586311513 wute = -5.1775069626344e-6   ua1 = 9.27458968906933e-09 wua1 = -1.12560876657858e-14   ub1 = -4.47182091258746e-18 wub1 = 5.86524560975631e-24   uc1 = 4.207051006468e-10 wuc1 = -4.87191718685898e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.55 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.22018585571533+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.5646314332372e-7   k1 = 0.214861425044933 wk1 = 3.27040736184641e-7   k2 = 0.0520850050141133 wk2 = -4.94706122707028e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 47987.59018134 wvsat = 0.00856282383240925   ua = 3.44169001577159e-09 wua = -5.70494892075117e-15   ub = -1.64199871850573e-18 wub = 3.19923630495839e-24   uc = -2.7937238741136e-10 wuc = 2.83988436891214e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0260855438916973 wu0 = -2.50351605670567e-8   a0 = 0.783374013593333 wa0 = 5.86437040018102e-7   keta = -0.0200886954067375 wketa = 3.15679974876173e-8   a1 = 0.0   a2 = 0.8   ags = -0.0656680853125332 wags = 3.33227815138276e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.319878220519267+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.70274173315858e-7   nfactor = {2.43585188798533+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.15094816761619e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.594026026461021 wpclm = -6.99514514884491e-7   pdiblc1 = 0.39   pdiblc2 = -0.000946599370666533 wpdiblc2 = 1.78861484556857e-9   pdiblcb = 0.580662666666667 wpdiblcb = -9.51521608297866e-7   drout = 0.56   pscbe1 = 627343825.1902 wpscbe1 = 203.896855410189   pscbe2 = 7.15160495793333e-09 wpscbe2 = 4.2758050751277e-15   pvag = 0.0   delta = 0.01   alpha0 = 7.17677495617133e-11 walpha0 = -8.47607408314149e-17   alpha1 = 2.5401143235454e-16 walpha1 = -2.99998220893157e-22   beta0 = -51.856518105586 wbeta0 = 9.66760022277611e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -4.14462774745334e-11 wagidl = 2.22218070945401e-16   bgidl = 2420143596.69 wbgidl = -1677.24951775067   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.137583350960667 wkt1 = -4.81896691240042e-7   kt2 = -0.05321158589764 wkt2 = 8.59309649237788e-10   at = 332265.066666667 wat = -0.380608643319147   ute = 3.12434586311513 wute = -5.17750696263439e-6   ua1 = 9.27458968906933e-09 wua1 = -1.12560876657858e-14   ub1 = -4.47182091258746e-18 wub1 = 5.86524560975631e-24   uc1 = 4.207051006468e-10 wuc1 = -4.87191718685898e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.56 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.29508256927302+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.03865088805347e-07 wvth0 = 3.70186364364353e-07 pvth0 = -9.16909163444622e-13   k1 = -0.0469712570197247 lk1 = 2.11106213205643e-06 wk1 = 6.86670508393115e-07 pk1 = -2.89956466733939e-12   k2 = 0.121607739862363 lk2 = -5.60536643851424e-07 wk2 = -1.36904793072537e-07 pk2 = 7.04950148631738e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 106187.186466784 lvsat = -0.469242276595683 wvsat = -0.0451886861901439 pvsat = 4.33378967265218e-7   ua = 5.74737344679617e-09 lua = -1.85898908469492e-14 wua = -9.17512980429135e-15 pua = 2.79788122585046e-20   ub = -3.71794396203174e-18 lub = 1.6737595006372e-23 wub = 6.19352079492536e-24 pub = -2.41418319116183e-29   uc = -3.82229339039872e-10 luc = 8.29298366764206e-16 wuc = 4.24244415292864e-16 puc = -1.13083318118832e-21   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.031946398429509 lu0 = -4.7253948509033e-08 wu0 = -3.4608835136346e-08 pu0 = 7.7189072381985e-14   a0 = 0.720421733770763 la0 = 5.07561443484084e-07 wa0 = 7.33154390015627e-07 pa0 = -1.18292888134936e-12   keta = 0.00906378945981384 lketa = -2.35045932279482e-07 wketa = 1.23751324143653e-09 pketa = 2.44543714841658e-13   a1 = 0.0   a2 = 0.8   ags = -0.631668939101425 lags = 4.56345999179076e-06 wags = 9.47195010417289e-07 pags = -4.95019523940999e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.310601329247027+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.47962160934256e-08 wvoff = 1.61124863327408e-07 pvoff = 7.37675743866607e-14   nfactor = {6.10720753200998+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.96008115270276e-05 wnfactor = -6.84026410413934e-06 pnfactor = 4.58708948638172e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.374340329800135 lpclm = 7.80758738191273e-06 wpclm = 4.00667737133301e-07 ppclm = -8.87037123204423e-12   pdiblc1 = 0.39   pdiblc2 = 0.000404591556747858 lpdiblc2 = -1.08941633166265e-08 wpdiblc2 = -3.71038453002076e-10 ppdiblc2 = 1.7412502751881e-14   pdiblcb = 0.580662666666667 wpdiblcb = -9.51521608297866e-7   drout = 0.56   pscbe1 = 451983879.496263 lpscbe1 = 1413.86376182989 wpscbe1 = 410.986730269869 ppscbe1 = -0.00166969069445891   pscbe2 = 4.72933450123451e-09 lpscbe2 = 1.95298898304573e-14 wpscbe2 = 8.65892973302734e-15 ppscbe2 = -3.53395474255184e-20   pvag = 0.0   delta = 0.01   alpha0 = 8.50868922531286e-11 lalpha0 = -1.07387425991227e-16 walpha0 = -1.00491210417798e-16 palpha0 = 1.26829081845016e-22   alpha1 = -3.62202609688672e-12 lalpha1 = 2.92051332479775e-17 walpha1 = 4.2777656699245e-18 palpha1 = -3.44924948224845e-23   beta0 = -24.5272112950764 lbeta0 = -0.000220346307604073 wbeta0 = 6.43989375878019e-05 pbeta0 = 2.60238287894591e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.54539697142822e-10 lagidl = 9.11831302967491e-16 wagidl = 3.42866381831422e-16 pagidl = -9.72743655985441e-22   bgidl = 3862525932.03237 lbgidl = -11629.4066274601 wbgidl = -3380.76392432456 pbgidl = 0.0137348199879901   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.156764145155264 lkt1 = -2.37321730738915e-06 wkt1 = -9.30690438086097e-07 pkt1 = 3.61846151748338e-12   kt2 = 0.0209028649696082 lkt2 = -5.97557987911408e-07 wkt2 = -1.17551458966987e-07 pkt2 = 9.54703162654381e-13   at = 650204.028482641 lat = -2.56342675521802 wat = -0.810409202724985 pat = 3.46532632268677e-6   ute = 6.71890076326217 lute = -2.89815949310117e-05 wute = -1.08496769306534e-05 pute = 4.57326531266091e-11   ua1 = 1.56738625512061e-08 lua1 = -5.15950205506325e-14 wua1 = -2.14236710526285e-14 pua1 = 8.19775441829267e-20   ub1 = -8.35994043663327e-18 lub1 = 3.13485002231136e-23 wub1 = 1.22683873832211e-23 pub1 = -5.16262141821248e-29   uc1 = 1.1352187167731e-09 luc1 = -5.76086463289729e-15 wuc1 = -1.22526918992045e-15 puc1 = 5.95085146651959e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.57 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.20077550984404+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.20729645500891e-07 wvth0 = 2.17497806022171e-07 pvth0 = -2.96590824158454e-13   k1 = 0.26854496287297 lk1 = 8.29233947504013e-07 wk1 = 2.00040806572495e-07 pk1 = -9.2256434879427e-13   k2 = 0.0713502107333985 lk2 = -3.56358496225985e-07 wk2 = -6.6892138681257e-08 pk2 = 4.20514078420857e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 45714.7670748441 lvsat = -0.22356472762205 wvsat = -0.016529372207623 pvsat = 3.16946549225897e-7   ua = 2.49808158056208e-09 lua = -5.38919423809566e-15 wua = -3.54401405534183e-15 pua = 5.10162743442384e-21   ub = -4.34508992764776e-19 lub = 3.39818732969923e-24 wub = 1.06229582772575e-24 pub = -3.29552237332444e-30   uc = -2.34424038354754e-10 luc = 2.28818935599417e-16 wuc = 2.0079656102345e-16 puc = -2.2304543741494e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0258290445612361 lu0 = -2.24013542243405e-08 wu0 = -2.08329175006763e-08 pu0 = 2.12225059104432e-14   a0 = 1.08433562796474 la0 = -9.70888971796338e-07 wa0 = 2.67049701325564e-07 pa0 = 7.10685738901055e-13   keta = -0.0236350473119817 lketa = -1.02202395454588e-07 wketa = 4.15086198144555e-08 pketa = 8.09367869760613e-14   a1 = 0.0   a2 = 0.8   ags = -0.0391856616103867 lags = 2.15641491429112e-06 wags = 2.13328638402491e-07 pags = -1.96876182954054e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.408879048410286+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.24470580332558e-07 wvoff = 2.81400290617226e-07 pvoff = -4.14867946987195e-13   nfactor = {-3.92690538510466+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.11641569063332e-05 wnfactor = 8.9050020465192e-06 pnfactor = -1.8096421719962e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.16829098775029 leta0 = 1.00871640189186e-06 weta0 = 3.90075619635389e-07 peta0 = -1.58473603520428e-12   etab = 0.147059412310586 letab = -8.81833816710654e-07 wetab = -3.4100949664713e-07 petab = 1.3853981394395e-12   dsub = -0.376947123586 ldsub = 3.80647698827118e-06 wdsub = 1.47198347032222e-06 pdsub = -5.98013598190293e-12   voffl = 0.0   minv = 0.0   pclm = 2.51628487330623 lpclm = -3.93597641198492e-06 wpclm = -3.30976221533642e-06 ppclm = 6.20376248919745e-12   pdiblc1 = 0.39   pdiblc2 = -0.00484696072685175 lpdiblc2 = 1.0440992549712e-08 wpdiblc2 = 7.95255391662678e-09 ppdiblc2 = -1.64032399054832e-14   pdiblcb = 0.482358059867636 lpdiblcb = 3.99376031156801e-07 wpdiblcb = -8.35419719213804e-07 ppdiblcb = -4.71679946464697e-13   drout = 0.56   pscbe1 = 800000123.029408 lpscbe1 = -0.000253765132583794 wpscbe1 = -0.000193284392480564 ppscbe1 = 3.986757313168e-10   pscbe2 = 1.11138847422396e-08 lpscbe2 = -6.40822659155922e-15 wpscbe2 = -1.74341102455455e-15 ppscbe2 = 6.92139742518247e-21   pvag = 0.0   delta = 0.01   alpha0 = -8.0854915868073e-11 lalpha0 = 5.66774069470676e-16 walpha0 = 9.17793062382925e-17 palpha0 = -6.5429642540165e-22   alpha1 = -4.08211663342731e-10 lalpha1 = 1.67290636792916e-15 walpha1 = 4.82118762293449e-16 palpha1 = -1.97578748566309e-21   beta0 = -177.700038792644 lbeta0 = 0.000401939441954988 wbeta0 = 0.000278189354793618 pbeta0 = -6.0831478508161e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.57534074211767e-10 lagidl = -7.62275259340974e-16 wagidl = -2.28893504570667e-16 pagidl = 1.35010978538737e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.367244975244181 lkt1 = -2.44357942507792e-07 wkt1 = -9.92566095988537e-08 pkt1 = 2.40646851385622e-13   kt2 = -0.165027115726472 lkt2 = 1.57808217003753e-07 wkt2 = 1.862037105989e-07 pkt2 = -2.79344131920436e-13   at = -50754.1561642239 lat = 0.284312602139347 wat = 0.183450087627019 pat = -5.72364196950313e-7   ute = 0.712203472727261 lute = -4.57855826398756e-06 wute = 8.11213813315737e-08 pute = 1.32477653400296e-12   ua1 = 6.2929410245608e-09 lua1 = -1.34837322814654e-14 wua1 = -2.64023112445909e-15 pua1 = 5.66722736002852e-21   ub1 = -1.52914047797682e-18 lub1 = 3.59743274067747e-24 wub1 = -1.53977142710682e-24 pub1 = 4.47133651074832e-30   uc1 = -4.2319640390823e-10 luc1 = 5.70411856157249e-16 wuc1 = 2.32532213078817e-16 puc1 = 2.83320902414617e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.58 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.14901642035076+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.13969380666659e-07 wvth0 = 1.29520817061055e-07 pvth0 = -1.15126143601672e-13   k1 = 0.784819192725983 lk1 = -2.35652897411546e-07 wk1 = -3.7259505643399e-07 pk1 = 2.58576142405701e-13   k2 = -0.193119342046643 lk2 = 1.89146453181134e-07 wk2 = 2.54016268529233e-07 pk2 = -2.41403796810973e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -343848.453230798 lvsat = 0.579963173982739 wvsat = 0.500118684728169 pvsat = -7.48711365636032e-7   ua = 3.1342242540839e-09 lua = -6.70132628992338e-15 wua = -5.27169039253842e-15 pua = 8.66519829922634e-21   ub = -6.81657926646484e-19 lub = 3.90796611238313e-24 wub = 1.90867795606258e-24 pub = -5.04130231375284e-30   uc = -2.82529724407897e-10 luc = 3.28043551668701e-16 wuc = 2.85071981281946e-16 puc = -3.96875121706084e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0287146507375326 lu0 = -2.83533151766044e-08 wu0 = -2.84811778910427e-08 pu0 = 3.69980984255077e-14   a0 = -1.36726104114786 la0 = 4.08586747858875e-06 wa0 = 3.48673753987238e-06 pa0 = -5.93036474502348e-12   keta = -0.238858055470237 lketa = 3.41724759646939e-07 wketa = 3.17864584587657e-07 pketa = -4.89085527491805e-13   a1 = 0.0   a2 = 0.8   ags = 3.12984028065267 lags = -4.38013841720648e-06 wags = -4.13651939059229e-06 pags = 7.0034000092892e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.285177019718355+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.93180752754917e-08 wvoff = 1.38632071874224e-07 pvoff = -1.20388793815567e-13   nfactor = {3.49163218630427+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.13760059288256e-06 wnfactor = -2.68132423175869e-06 pnfactor = 5.80197514201257e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -1.17847994230115 leta0 = 3.09237052672875e-06 weta0 = 1.292650949266e-06 peta0 = -3.4464222079629e-12   etab = 96.8844326556782 letab = -0.000200416015888664 wetab = -0.000114417036382055 petab = 2.36682946082304e-10   dsub = 3.718085894344 ldsub = -4.64009372576592e-06 wdsub = -4.46065146884209e-06 pdsub = 6.25674228374506e-12   voffl = 0.0   minv = 0.0   pclm = -0.234685206685917 lpclm = 1.73827901186993e-06 wpclm = 6.69282295956371e-07 ppclm = -2.00356592348649e-12   pdiblc1 = 0.424522071657199 lpdiblc1 = -7.12065368388627e-08 wpdiblc1 = -3.10322249014898e-08 ppdiblc1 = 6.40082463063587e-14   pdiblc2 = -0.000705337347139934 lpdiblc2 = 1.89832278503002e-09 wpdiblc2 = 1.08695724520831e-09 ppdiblc2 = -2.24199931834198e-15   pdiblcb = 1.31718254415305 lpdiblcb = -1.32256467346071e-06 wpdiblcb = -2.07238672901284e-06 ppdiblcb = 2.07973521269317e-12   drout = 0.836726016187682 ldrout = -5.7078559657733e-07 wdrout = -7.67654504877351e-07 pdrout = 1.58339335263121e-12   pscbe1 = 800000000.0   pscbe2 = 1.20412358400074e-08 lpscbe2 = -8.32101620515684e-15 wpscbe2 = -1.94464758375744e-15 ppscbe2 = 7.33647559918359e-21   pvag = 0.0   delta = 0.01   alpha0 = 2.93735847514385e-10 lalpha0 = -2.05871073530991e-16 walpha0 = -4.64988940740911e-16 palpha0 = 4.9411491801104e-22   alpha1 = 7.24649679075235e-10 lalpha1 = -6.6377648567315e-16 walpha1 = -9.81351006043651e-16 palpha1 = 1.04282087036021e-21   beta0 = 26.0525115679886 lbeta0 = -1.83283110157657e-05 wbeta0 = -3.46318967754458e-05 pbeta0 = 3.69222156123001e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -3.37339491576963e-10 lagidl = 4.64733562650361e-16 wagidl = 8.77985344906736e-16 pagidl = -9.32980590941005e-22   bgidl = 150624086.835614 lbgidl = 1751.95503477756 wbgidl = 1003.14879711067 pbgidl = -0.00206913282857477   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.730878175417046 lkt1 = 5.05685714230368e-07 wkt1 = 3.6077369075444e-07 pkt1 = -7.08229127274495e-13   kt2 = -0.173267439165446 lkt2 = 1.74805021261273e-07 wkt2 = 1.73889604589859e-07 pkt2 = -2.5394458893016e-13   at = -23876.965133592 lat = 0.228874686586306 wat = 0.0175687188778979 pat = -2.30210982276364e-7   ute = -5.20842596217808 lute = 7.63355699236674e-06 wute = 5.46875388180494e-06 pute = -9.78795899150842e-12   ua1 = -2.35692998253048e-09 lua1 = 4.35782035285937e-15 wua1 = 2.71194626283449e-15 pua1 = -5.37237710174395e-21   ub1 = -2.0616127911522e-19 lub1 = 8.68605571895976e-25 wub1 = 1.46015961818302e-24 pub1 = -1.71643526064623e-30   uc1 = -5.54187330662127e-10 luc1 = 8.40598719335054e-16 wuc1 = 7.4569420130752e-16 puc1 = -1.03013532683461e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.59 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05799279108544+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.72442133114233e-08 wvth0 = 7.8125552835867e-09 pvth0 = 1.42056802770154e-14   k1 = 0.888609729582197 lk1 = -3.4594466591536e-07 wk1 = -5.8751690941158e-07 pk1 = 4.86960270410102e-13   k2 = -0.120647075196019 lk2 = 1.12134668479521e-07 wk2 = 1.70709389722211e-07 pk2 = -1.52878741729237e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 421449.457653882 lvsat = -0.233271467443935 wvsat = -0.525795690199018 pvsat = 3.41464233907845e-7   ua = -5.1755448160878e-09 lua = 2.12895009526575e-15 wua = 5.78154680244987e-15 pua = -3.08039156718163e-21   ub = 4.55576487131242e-18 lub = -1.65751837479433e-24 wub = -5.12925395871218e-24 pub = 2.43747158029958e-30   uc = 1.37970483617899e-11 luc = 1.31554625062659e-17 wuc = -1.09514884958001e-16 puc = 2.2427876661401e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00393713159004925 lu0 = 6.34370949241257e-09 wu0 = 1.48905978429207e-08 pu0 = -9.09039859687963e-15   a0 = 4.57859399163621 la0 = -2.23242402173887e-06 wa0 = -5.14749148173078e-06 pa0 = 3.24469511403486e-12   keta = 0.1183345492966 lketa = -3.78416754972835e-08 wketa = -1.90408862116119e-07 pketa = 5.10251513666017e-14   a1 = 0.0   a2 = 0.613277635331865 la2 = 1.98418280146217e-07 wa2 = 2.20526992356855e-07 pa2 = -2.34340362104105e-13   ags = -2.17998841309484 lags = 1.26228732626e-06 wags = 3.55545315498465e-06 pags = -1.17038231259759e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.22274284177294+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.97314529193086e-09 wvoff = 1.39443411466191e-08 pvoff = 1.21091269893542e-14   nfactor = {-1.1937174323113+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.41229955143849e-07 wnfactor = 3.77974549811651e-06 pnfactor = -1.06380307360256e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 3.12876067560346 leta0 = -1.48466702900018e-06 weta0 = -4.14560437707356e-06 peta0 = 2.33247455550791e-12   etab = -194.923781655119 letab = 0.000109670481350133 wetab = 0.000230195649940023 petab = -1.29515589685617e-10   dsub = -1.60807359420033 ldsub = 1.01968574082185e-06 wdsub = 2.88297686975126e-06 pdsub = -1.54687624672109e-12   voffl = 0.0   minv = 0.0   pclm = 2.28844924895913 lpclm = -9.42899539807812e-07 wpclm = -2.60283970653907e-06 ppclm = 1.47351525700126e-12   pdiblc1 = 0.431214614239296 lpdiblc1 = -7.83182869032164e-08 wpdiblc1 = 2.43957295620762e-07 ppdiblc1 = -2.28206067802366e-13   pdiblc2 = 0.00144842800847288 lpdiblc2 = -3.90350124927667e-10 wpdiblc2 = -1.87827853493819e-09 ppdiblc2 = 9.08972900601333e-16   pdiblcb = 1.08897186468201 lpdiblcb = -1.08005933344896e-06 wpdiblcb = -1.31564778180215e-06 ppdiblcb = 1.27559565130709e-12   drout = -0.488573472375366 ldrout = 8.37528001350331e-07 wdrout = 1.5353090097547e-06 pdrout = -8.63823190630366e-13   pscbe1 = 800000000.0   pscbe2 = -1.56308948108599e-09 lpscbe2 = 6.13545684539924e-15 wpscbe2 = 1.057268260655e-14 ppscbe2 = -5.96491511958431e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.94276274285744 lbeta0 = 1.97843425627414e-06 wbeta0 = 2.13888157049548e-06 pbeta0 = -2.15181074767424e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.61020264673129e-10 lagidl = -4.89897652011725e-16 wagidl = -9.14431105571545e-16 pagidl = 9.71709241162336e-22   bgidl = 2698751826.32877 lbgidl = -955.782330061967 wbgidl = -2006.29759422135 pbgidl = 0.00112881926581751   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.030211418283097 lkt1 = -3.03077009439965e-07 wkt1 = -6.49714588157156e-07 pkt1 = 3.65554116451566e-13   kt2 = 0.043470644370762 lkt2 = -5.55091023514768e-08 wkt2 = -1.38325774576002e-07 pkt2 = 7.78273371558927e-14   at = 293608.56910877 lat = -0.108497506549929 wat = -0.37554342330991 pat = 1.87524918273803e-7   ute = 4.81758470563444 lute = -3.02046293165623e-06 wute = -8.36553551339007e-06 pute = 4.91288262282282e-12   ua1 = 3.08062421620629e-09 lua1 = -1.42033136577787e-15 wua1 = -4.98111989779605e-15 pua1 = 2.80256733705618e-21   ub1 = 1.28655772118657e-18 lub1 = -7.17614361146715e-25 wub1 = -1.04781673955123e-24 pub1 = 9.48635720183773e-31   uc1 = 4.76029692989825e-10 luc1 = -2.54149038244409e-16 wuc1 = -4.75464664291185e-16 puc1 = 2.67514487787464e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.60 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.12139301139888+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.29155864681326e-08 wvth0 = 1.31760133469284e-07 pvth0 = -5.55319372182309e-14   k1 = -1.06929827036745 lk1 = 7.55648775360312e-07 wk1 = 1.75911444312106e-06 pk1 = -8.33343700516155e-13   k2 = 0.569940425456 lk2 = -2.7641610171233e-07 wk2 = -6.54402790078942e-07 pk2 = 3.11360724889725e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 127862.754896356 lvsat = -0.0680884321778461 wvsat = -0.163037939946194 pvsat = 1.37362938821097e-7   ua = 4.56514718174584e-10 lua = -1.03986061697258e-15 wua = -1.22170871750098e-15 pua = 8.59906112052475e-22   ub = -1.78485319482925e-19 lub = 1.00615068405438e-24 wub = 6.65635298157114e-25 pub = -8.22953321406848e-31   uc = 1.16292433876398e-10 luc = -4.4512336208902e-17 wuc = -1.95364442595968e-16 puc = 7.07301000717113e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0101874331001463 lu0 = -1.60330733574966e-09 wu0 = -1.79584905079696e-09 pu0 = 2.98030510507868e-16   a0 = 1.92678787338843 la0 = -7.40417130980166e-07 wa0 = -4.57443594519694e-07 pa0 = 6.05895950870192e-13   keta = 0.465517757121073 lketa = -2.33180141181229e-07 wketa = -6.23733440487353e-07 pketa = 2.94830025492236e-13   a1 = 0.0   a2 = 0.127167227846878 la2 = 4.71922467592756e-07 wa2 = 1.20269212303668e-06 pa2 = -7.86943786899542e-13   ags = -2.8166562312453 lags = 1.62050083412853e-06 wags = 6.1926640776134e-06 pags = -2.65417739168358e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.149650848646917+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.81511875365084e-08 wvoff = -6.20288634019902e-08 pvoff = 5.48545388501748e-14   nfactor = {-2.08445705789424+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.34239391660259e-06 wnfactor = 4.80138344499013e-06 pnfactor = -1.63861540475563e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.4829665674717 leta0 = -5.58680723589144e-07 weta0 = -1.17273541937323e-06 peta0 = 6.59825510885314e-13   etab = -0.00416606100549866 letab = 1.29867149223224e-09 wetab = 4.99599104256616e-09 petab = -1.58052907046338e-15   dsub = 0.309702812129811 ldsub = -5.93281408829272e-08 wdsub = -4.49602730090839e-07 pdsub = 3.28159674174863e-13   voffl = 0.0   minv = 0.0   pclm = -0.485677482136969 lpclm = 6.17929575922637e-07 wpclm = 1.29706838901419e-06 ppclm = -7.20721234064638e-13   pdiblc1 = 0.456130702636144 lpdiblc1 = -9.23370250466425e-08 wpdiblc1 = -8.08596680808352e-07 ppdiblc1 = 3.64000796387758e-13   pdiblc2 = 0.00447486484823391 lpdiblc2 = -2.09313849557715e-09 wpdiblc2 = -2.02165373826696e-08 ppdiblc2 = 1.12267741821712e-14   pdiblcb = -2.09306880417521 lpdiblcb = 7.10277664395533e-07 wpdiblcb = 2.73786746729334e-06 ppdiblcb = -1.0050660614135e-12   drout = 0.933750979925874 ldrout = 3.72742161564662e-08 wdrout = 9.17626380714124e-07 pdrout = -5.16291471592233e-13   pscbe1 = 799730588.317148 lpscbe1 = 0.151581250415802 wpscbe1 = 0.423257122931318 ppscbe1 = -2.38140541131745e-7   pscbe2 = 9.42200213820054e-09 lpscbe2 = -4.51731330928997e-17 wpscbe2 = 3.49081413833378e-17 ppscbe2 = -3.59627700518693e-23   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 13.7838779043953 lbeta0 = -1.87063709598319e-06 wbeta0 = -5.9982016333581e-06 pbeta0 = 2.42642147197554e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.32291358873614e-08 lagidl = 7.26896822505668e-15 wagidl = 1.64821654083831e-14 pagidl = -8.81627702825607e-21   bgidl = 2050367757.07247 lbgidl = -590.976814103738 wbgidl = -1650.17207188019 pbgidl = 0.000928449514178528   cgidl = 1505.10589248037 lcgidl = -0.00067803836913337 wcgidl = -0.00142328091448798 pcgidl = 8.00791927165688e-10   egidl = -6.27702854070459 legidl = 3.58795858408495e-06 wegidl = 7.53153981717654e-06 pegidl = -4.23753049965658e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.392513456940738 lkt1 = -6.5235931093777e-08 wkt1 = -1.31605953883192e-07 pkt1 = 7.40465106809318e-14   kt2 = 0.115733559927401 lkt2 = -9.6166964634433e-08 wkt2 = -2.57393163512417e-07 pkt2 = 1.448191747323e-13   at = 195683.792777014 lat = -0.0534013062441824 wat = -0.156641215616027 pat = 6.43622179413325e-8   ute = -0.429971460282673 lute = -6.79884255769576e-08 wute = 1.41856043425562e-07 pute = 1.26300852079184e-13   ua1 = 1.75897833029566e-09 lua1 = -6.76723167820893e-16 wua1 = -1.19355652841353e-15 pua1 = 6.71540258033531e-22   ub1 = -2.9074313186747e-19 lub1 = 1.69835036213903e-25 wub1 = 1.16090866346012e-24 pub1 = -2.94077123115726e-31   uc1 = 5.38760763423599e-11 luc1 = -1.66293716811127e-17 wuc1 = 1.67244275029693e-19 puc1 = -9.40979844141484e-26   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.61 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.746874846063829+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.41730237058862e-08 wvth0 = -4.07276811052895e-07 pvth0 = 1.12991495043295e-13   k1 = 3.37740378517193 lk1 = -6.34559261879408e-07 wk1 = -5.54862703076964e-06 pk1 = 1.45133397839809e-12   k2 = -1.01882103388497 lk2 = 2.20291103413111e-07 wk2 = 1.98431753001798e-06 pk2 = -5.13603518544737e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 89851.4690099752 lvsat = -0.0562046597808998 wvsat = -0.0900434406066304 pvsat = 1.14542084536574e-7   ua = -8.1132936247372e-09 lua = 1.63938712373868e-15 wua = 1.16059199008403e-14 pua = -3.1504980439285e-21   ub = 7.58306786078106e-18 lub = -1.42040577911699e-24 wub = -1.05125812984014e-23 pub = 2.67178195890802e-30   uc = -1.17616860759013e-10 luc = 2.86165978473236e-17 wuc = 1.38264822149083e-16 puc = -3.35750859996519e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00547556868789133 lu0 = 3.29354221725885e-09 wu0 = 2.04691967364576e-08 pu0 = -6.66286887432782e-15   a0 = -3.00122212343589 la0 = 8.00266058406996e-07 wa0 = 3.37836258846361e-06 pa0 = -5.93322822565345e-13   keta = -1.30096884157891 lketa = 3.19090696063137e-07 wketa = 1.37287552016917e-06 pketa = -3.293858067495e-13   a1 = 0.0   a2 = 5.13731966507317 la2 = -1.0944415700768e-06 wa2 = -6.11640005002578e-06 pa2 = 1.50128255190236e-12   ags = 6.23727947577809 lags = -1.21010351744384e-06 wags = -1.02587897112383e-05 pags = 2.48917221795544e-12   b0 = 0.0   b1 = 2.21205892491735e-23 lb1 = -6.9157367816831e-30 wb1 = -3.47523791993178e-29 pb1 = 1.08649143281163e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.389127346544133+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 3.67182658130814e-08 wvoff = 4.04580567316191e-07 pvoff = -9.10253003506961e-14   nfactor = {-7.20271580632193+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.94255609519352e-06 wnfactor = 1.53302144738108e-05 pnfactor = -4.93032807994408e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -1.68058593065764 leta0 = 4.30366002321018e-07 weta0 = 3.70421012137159e-06 peta0 = -8.64892989082064e-13   etab = 0.762787687875484 letab = -2.38480214650421e-07 wetab = -7.72035360968816e-07 petab = 2.41348998759671e-13   dsub = -0.429421519934689 ldsub = 1.71750212045055e-07 wdsub = 2.71653877049784e-06 pdsub = -6.6169647228618e-13   voffl = 0.0   minv = 0.0   pclm = 4.37888484253035 lpclm = -9.02917460136707e-07 wpclm = -4.35734993297256e-06 ppclm = 1.04706480128466e-12   pdiblc1 = -0.208384808075712 lpdiblc1 = 1.15415775191292e-07 wpdiblc1 = 2.0595748491845e-06 ppdiblc1 = -5.32698614406147e-13   pdiblc2 = -0.0418430563041281 lpdiblc2 = 1.2387603737655e-08 wpdiblc2 = 9.83206875890269e-08 ppdiblc2 = -2.583246675853e-14   pdiblcb = 0.0140728948446869 lpdiblcb = 5.15050978973499e-08 wpdiblcb = -8.96424571952594e-07 ppdiblcb = 1.31151733152275e-13   drout = 1.23660364312187 ldrout = -5.74090347598047e-08 wdrout = -3.27723707397901e-06 pdrout = 7.95182249156119e-13   pscbe1 = 800962184.581608 lpscbe1 = -0.233462542512825 wpscbe1 = -1.5116325818999 ppscbe1 = 3.66779506407247e-7   pscbe2 = 7.65598425804173e-09 lpscbe2 = 5.06951164924198e-16 wpscbe2 = 1.10354770270716e-15 ppscbe2 = -3.70060105225032e-22   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.31860878969437 lbeta0 = 1.50651709498681e-07 wbeta0 = 4.3821703602206e-06 pbeta0 = -8.18877267352924e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.15964942320844e-08 lagidl = -9.87160712422662e-15 wagidl = -4.90091108401483e-14 pagidl = 1.16587845955323e-20   bgidl = -2720311836.08139 lbgidl = 900.518912540695 wbgidl = 5844.76689164334 pbgidl = -0.00141475321349954   cgidl = -4003.94961600131 lcgidl = 0.00104430172692733 wcgidl = 0.00508314612317135 pcgidl = -1.23336440903405e-9   egidl = 22.8751019310878 legidl = -5.52610518235528e-06 wegidl = -2.68983564899162e-05 pegidl = 6.52656342200028e-12   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.03290239398564 lkt1 = 1.34973985406066e-07 wkt1 = 1.13098426556616e-06 pkt1 = -3.20687170347275e-13   kt2 = -0.413599271718949 lkt2 = 6.93225931858185e-08 wkt2 = 8.86938756259448e-07 pkt2 = -2.12942468001337e-13   at = -221994.135888449 lat = 0.0771806860179307 wat = 0.3711331029686 pat = -1.00640089472328e-7   ute = -0.971688022730622 lute = 1.01372757073644e-07 wute = 1.05525022894437e-06 pute = -1.59260879293044e-13   ua1 = -2.11136085673731e-09 lua1 = 5.33291934934723e-16 wua1 = 4.00082333262634e-15 pua1 = -9.52420272962253e-22   ub1 = 2.52489092666666e-19 wub1 = 2.20277252320957e-25   uc1 = 4.55904165152093e-12 luc1 = -1.21099258943818e-18 wuc1 = -6.21911453710708e-18 puc1 = 1.90252046189466e-24   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.62 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.82447466112572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.972936402211e-07 wvth0 = 1.3804446707427e-06 pvth0 = -3.20777669856622e-13   k1 = -3.45103748326211 lk1 = 1.02228007061089e-06 wk1 = 3.8467967691289e-06 pk1 = -8.28352861561697e-13   k2 = 1.69144245131634 lk2 = -4.37321808109164e-07 wk2 = -1.62629982671601e-06 pk2 = 3.62469455658485e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1542471.2433662 lvsat = 0.33985885850463 wvsat = 2.87971851809328 pvsat = -6.06035017598456e-7   ua = 7.51989918598393e-09 lua = -2.15381951346907e-15 wua = -1.27662531567666e-14 pua = 2.76311728242311e-21   ub = -6.10129214587244e-18 lub = 1.89993996417741e-24 wub = 9.98947684575904e-24 pub = -2.30279642507479e-30   uc = 3.4569726900288e-12 luc = -7.60514953085039e-19 wuc = -3.24462578439213e-18 puc = 7.60483428030604e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0296638344401482 lu0 = -5.23261227892241e-09 wu0 = -3.58989420094699e-08 pu0 = 7.01418357470654e-15   a0 = -1.10058616375073 la0 = 3.39099550420906e-07 wa0 = 4.04146028482904e-06 pa0 = -7.54215521416054e-13   keta = -1.11998101488211 lketa = 2.75176171769079e-07 wketa = 1.75314180010364e-06 pketa = -4.21652856380238e-13   a1 = 0.0   a2 = -4.71644684406887 la2 = 1.29645662816841e-06 wa2 = 4.81705494816764e-06 pa2 = -1.15158910194929e-12   ags = 1.25   b0 = 0.0   b1 = -5.16147082480718e-23 lb1 = 1.09752483324535e-29 wb1 = 8.10888847984088e-29 pb1 = -1.72425782857641e-35   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.01602494898349+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.88827446273763e-07 wvoff = 7.47209581620675e-07 pvoff = -1.74160119123508e-13   nfactor = {33.6689548729063+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -6.97446433507305e-06 wnfactor = -4.76950364469032e-05 pnfactor = 1.03619927529561e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -3.32030265215721 leta0 = 8.2822358819223e-07 weta0 = 4.1771021349569e-06 peta0 = -9.79634561474376e-13   etab = -1.0871077021341 letab = 2.10374702990724e-07 wetab = 1.10579788884361e-06 petab = -2.14284705308317e-13   dsub = 0.409011776371377 ldsub = -3.16855661040574e-08 wdsub = -8.53646030041823e-08 pdsub = 1.81517584536034e-14   voffl = 0.0   minv = 0.0   pclm = 4.84261104945823 lpclm = -1.01543505953327e-06 wpclm = -4.93645429098318e-06 ppclm = 1.18757752450364e-12   pdiblc1 = 4.65621739491621 lpdiblc1 = -1.06492157413826e-06 wpdiblc1 = -5.23490812208694e-06 ppdiblc1 = 1.23722014477721e-12   pdiblc2 = 0.119119015306646 lpdiblc2 = -2.666791139384e-08 wpdiblc2 = -1.40763507512405e-07 ppdiblc2 = 3.21784441724913e-14   pdiblcb = -1.4288416749563 lpdiblcb = 4.01611003284721e-07 wpdiblcb = 2.24258232792022e-06 ppdiblcb = -6.30490623019066e-13   drout = 1.0   pscbe1 = 800000000.0   pscbe2 = 9.65288895901301e-09 lpscbe2 = 2.24262020899211e-17 wpscbe2 = 1.44160786941811e-15 ppscbe2 = -4.52086347955425e-22   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 19.3830832798952 lbeta0 = -2.77664825185468e-06 wbeta0 = -5.35710966057581e-06 pbeta0 = 1.54424215833307e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.92373424114671e-09 lagidl = -1.70131598554548e-15 wagidl = -1.1758115174643e-14 pagidl = 2.62027750924541e-21   bgidl = 927662975.252689 lbgidl = 15.3816002682188 wbgidl = 113.64451850047 pbgidl = -2.41651431249022e-5   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 1.17581870713931 lkt1 = -4.00945685128689e-07 wkt1 = -1.54224700396111e-06 pkt1 = 3.27940318428284e-13   kt2 = -0.183858230184125 lkt2 = 1.35786863498919e-08 wkt2 = 7.54192646647647e-08 pkt2 = -1.60370015997864e-14   at = 750690.925009233 lat = -0.158829671788161 wat = -0.748085942724269 pat = 1.70924981336498e-7   ute = -2.97416636818895 lute = 5.87250097858963e-07 wute = 3.22609752525199e-06 pute = -6.85990925574533e-13   ua1 = -7.49432394937515e-11 lua1 = 3.91796371219803e-17 wua1 = -6.05547717172931e-18 pua1 = 1.98007876895318e-23   ub1 = -5.72694537118185e-19 lub1 = 2.00220905563736e-25 wub1 = 1.78158773162175e-24 pub1 = -3.78833252076585e-31   uc1 = -4.9199024013215e-11 luc1 = 1.1832756947322e-17 wuc1 = 1.31175649613359e-17 puc1 = -2.78929277824855e-24   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.63 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.003036+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.010197753   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.38874612e-9   ub = 1.066826e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0048880282   a0 = 1.279916   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21647917   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17570541+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4613328+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.64 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.003036+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.010197753   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.38874612e-9   ub = 1.066826e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0048880282   a0 = 1.279916   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21647917   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17570541+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4613328+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.65 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.981642148292+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.72490881747276e-7   k1 = 0.534439388927655 lk1 = -3.44027675352128e-7   k2 = 0.005689110475084 lk2 = 3.63515525498037e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 67925.4832099965 lvsat = -0.102296059716034   ua = -2.02129883628681e-09 lua = 5.10004356733726e-15   ub = 1.52617076555832e-18 lub = -3.7035305618916e-24   uc = -2.30174367955125e-11 luc = -1.28189165170151e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0026427586981379 lu0 = 1.81027952059545e-8   a0 = 1.341190737635 la0 = -4.94036028095979e-7   keta = 0.0101116040437775 lketa = -2.79883734203168e-8   a1 = 0.0   a2 = 0.8   ags = 0.170330354757245 lags = 3.72081191431215e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.174175329119845+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.23364882474108e-8   nfactor = {0.315488909136601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.2385244965431e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.0350910319060362 lpclm = 2.96957167307167e-07 wpclm = 4.96308367531817e-24 ppclm = -7.57306469012171e-29   pdiblc1 = 0.39   pdiblc2 = 9.04296639703799e-05 lpdiblc2 = 3.8491733328861e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799970369.961946 lpscbe1 = 0.120294865781034   pscbe2 = 1.20609351273826e-08 lpscbe2 = -1.03924511540718e-14   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.35768627006325e-10 lagidl = 8.81997206366977e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.631260565634999 lkt1 = 6.90569505210245e-7   kt2 = -0.078629106849 lkt2 = 2.10798531994808e-7   at = -35977.38207575 lat = 0.370698987864461 wat = 1.38777878078145e-17   ute = -2.46762697525 lute = 9.7406904594757e-6   ua1 = -2.465769591175e-09 lua1 = 1.7816169145152e-14 pua1 = -3.00926553810506e-36   ub1 = 2.02782333948e-18 lub1 = -1.23639210452584e-23 wub1 = 7.3468396926393e-40   uc1 = 9.777129116845e-11 luc1 = -7.22220402810009e-16 wuc1 = 1.23259516440783e-32 puc1 = -9.4039548065783e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.66 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0166179869188+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.03967106601765e-8   k1 = 0.43792147335879 lk1 = 4.8089676118731e-8   k2 = 0.01471198164958 lk2 = -3.05106752808383e-10   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 31719.18570813 lvsat = 0.0447970203543543   ua = -5.02669836569194e-10 lua = -1.06959631481753e-15   ub = 4.6494729061422e-19 lub = 6.07836253908346e-25   uc = -6.4407623172087e-11 luc = 3.99641788304033e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00818960923819999 lu0 = -4.43205057842235e-9   a0 = 1.3104492260441 la0 = -3.69144394929349e-7   keta = 0.0115107076952954 lketa = -3.36724250809121e-08 pketa = -6.31088724176809e-30   a1 = 0.0   a2 = 0.8   ags = 0.14144178625091 lags = 4.89444987610655e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17061466580209+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.68021743473288e-8   nfactor = {3.6130470793536+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.15826063299095e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.1619898605 leta0 = -3.33095122881999e-7   etab = -0.141676668963335 letab = 2.91196359043864e-7   dsub = 0.869395700000001 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = -0.286123216206924 lpclm = 1.31681005847096e-06 wpclm = -5.29395592033938e-23 ppclm = 2.01948391736579e-28   pdiblc1 = 0.39   pdiblc2 = 0.0018865445760297 lpdiblc2 = -3.44779136121275e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799999959.37362 lpscbe1 = 8.37975148897385e-5   pscbe2 = 9.6377215496335e-09 lpscbe2 = -5.4781159099233e-16   pvag = 0.0   delta = 0.01   alpha0 = -3.144478223853e-12 lalpha0 = 1.27748767223977e-17   alpha1 = 3.0154328869995e-15 lalpha1 = -1.22506122331739e-20   beta0 = 57.845613 lbeta0 = -0.000113126645507094   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37277016954699e-11 lagidl = 3.8087592135974e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.45128651889 lkt1 = -4.05998961097667e-8   kt2 = -0.007366609947 lkt2 = -7.87151958941399e-8   at = 104574.830071 lat = -0.200313770186987   ute = 0.78088974095 lute = -3.45685699539363e-06 wute = -2.11758236813575e-22 pute = -6.05845175209737e-28   ua1 = 4.05743146829e-09 lua1 = -8.68523536067074e-15   ub1 = -2.83288002861e-18 lub1 = 7.38335716467207e-24 wub1 = 1.46936793852786e-39 pub1 = -2.80259692864963e-45   uc1 = -2.26309101254e-10 luc1 = 5.94400914500348e-16 wuc1 = -9.86076131526265e-32   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.67 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0393498757844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.64909471257819e-8   k1 = 0.46933930857452 lk1 = -1.67139446749717e-8   k2 = 0.021958720811088 lk2 = -1.52525063234229e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 79606.936194042 lvsat = -0.0539780735324064 wvsat = 5.55111512312578e-17   ua = -1.32936764173355e-09 lua = 6.35581992631081e-16   ub = 9.3443839579024e-19 lub = -3.60553940289708e-25 wub = 7.3468396926393e-40   uc = -4.1156485346714e-11 luc = -7.99450159144852e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00459935842110001 lu0 = 2.97333718645914e-9   a0 = 1.5849937892658 la0 = -9.3543044372383e-7   keta = 0.0302810020398646 lketa = -7.23887474672056e-08 wketa = -6.61744490042422e-24 pketa = 6.31088724176809e-30   a1 = 0.0   a2 = 0.8   ags = -0.37259120790234 lags = 1.54970897460493e-06 pags = -4.03896783473158e-28   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1677958864496+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.26162957533899e-8   nfactor = {1.2213286935428+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.74988594881067e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.083979721 leta0 = 1.74251082763998e-07 weta0 = 1.65436122510606e-23 peta0 = -3.31321580192825e-29   etab = 0.00640714392666938 letab = -1.42469406079481e-08 wetab = -8.27180612553028e-25 petab = 5.52202633654708e-30   dsub = -0.0587913999999996 ldsub = 6.575512557132e-7   voffl = 0.0   minv = 0.0   pclm = 0.33200266945972 lpclm = 4.1840117911282e-8   pdiblc1 = 0.39824678284746 lpdiblc1 = -1.70101276789198e-8   pdiblc2 = 0.000215   pdiblcb = -0.4375276 lpdiblcb = 4.383675038088e-7   drout = 0.1867454271136 ldrout = 7.69889065709258e-7   pscbe1 = 800000000.0   pscbe2 = 1.039468368145e-08 lpscbe2 = -2.10915044863808e-15   pvag = 0.0   delta = 0.01   alpha0 = -9.9974843552294e-11 lalpha0 = 2.12500867802723e-16 walpha0 = 2.1570415377137e-32 palpha0 = -6.46521892952258e-38   alpha1 = -1.06269830865774e-10 lalpha1 = 2.19190160531544e-16 walpha1 = -2.18171751512617e-32 palpha1 = 8.18483859508097e-38   beta0 = -3.2706546791156 lbeta0 = 1.29340906260216e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.0605930052948e-10 lagidl = -3.25230242996046e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.42540755738626 lkt1 = -9.39788255079182e-8   kt2 = -0.02603340757042 lkt2 = -4.02123497777641e-8   at = -9001.358759918 lat = 0.0339527927908398   ute = -0.577978479603001 lute = -6.54003766688627e-7   ua1 = -6.06985160896602e-11 lua1 = -1.91023965949856e-16   ub1 = 1.03017017304036e-18 lub1 = -5.84716977159624e-25 wub1 = -7.3468396926393e-40   uc1 = 7.7199254260512e-11 luc1 = -3.16269529013939e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.68 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05137782399656+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.9272301958057e-8   k1 = 0.39115340718188 lk1 = 6.63693652091012e-8   k2 = 0.0238942373178024 lk2 = -1.73092597130849e-08 wk2 = 1.32348898008484e-23 pk2 = -6.31088724176809e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -23746.903830084 lvsat = 0.0558496443231508   ua = -2.8025250354396e-10 lua = -4.79247619584433e-16   ub = 2.1277529929528e-19 lub = 4.06312689243503e-25   uc = -7.8930277518692e-11 luc = 3.21453653745979e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.008670883468956 lu0 = -1.35322004734447e-9   a0 = 0.220162530228 la0 = 5.14891115717578e-7   keta = -0.0428864994653479 lketa = 5.36181999729047e-9   a1 = 0.0   a2 = 0.8   ags = 0.830448601759201 lags = 2.71313157345808e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21093603152804+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.32260617324734e-8   nfactor = {2.00663010659672+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.95025280837248e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.38136316 leta0 = 4.9026202561608e-07 weta0 = 1.05879118406788e-22 peta0 = 1.0097419586829e-28   etab = -0.014869899025 letab = 8.36285376012795e-9   dsub = 0.83297116249952 ldsub = -2.90069530176165e-7   voffl = 0.0   minv = 0.0   pclm = 0.0845993725202803 lpclm = 3.04740262564414e-7   pdiblc1 = 0.63777564619968 lpdiblc1 = -2.71542599973796e-7   pdiblc2 = -0.000141928826311 lpdiblc2 = 3.79286134133468e-10   pdiblcb = -0.025   drout = 0.8113877057728 ldrout = 1.06120443999403e-7   pscbe1 = 800000000.0   pscbe2 = 7.38890444982521e-09 lpscbe2 = 1.08490478249725e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.75377472066438 lbeta0 = 1.56475017498219e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.132375100038e-10 lagidl = 3.32858081155418e-16 pagidl = 9.4039548065783e-38   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.51990828798748 lkt1 = 6.44124185670019e-9   kt2 = -0.0736511439751599 lkt2 = 1.03880663998961e-8   at = -24367.726158164 lat = 0.050281678710177   ute = -2.265596160714 lute = 1.1393229107318e-6   ua1 = -1.13693879534068e-09 lua1 = 9.5262985191289e-16 wua1 = 3.94430452610506e-31 pua1 = -1.88079096131566e-37   ub1 = 3.9936102359928e-19 lub1 = 8.56047957841485e-26   uc1 = 7.3449104174976e-11 luc1 = -2.76419009148001e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.69 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.00983041569376+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.8961512453858e-9   k1 = 0.420161160566559 lk1 = 5.00485008602519e-8   k2 = 0.0158511726935312 lk2 = -1.27839259190142e-08 pk2 = 3.15544362088405e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -10183.0659440801 lvsat = 0.0482181137026453   ua = -5.779180205548e-10 lua = -3.11769688424489e-16   ub = 3.85114607900801e-19 lub = 3.0934804532831e-25   uc = -4.91245534217428e-11 luc = 1.53755323801385e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00866687011704799 lu0 = -1.35096198305365e-9   a0 = 1.53946590088 la0 = -2.27399094139321e-7   keta = -0.0626034569112048 lketa = 1.64553295007124e-8   a1 = 0.0   a2 = 1.14549842976048 la2 = -1.94390545523577e-07 wa2 = 8.470329472543e-22   ags = 2.42673310540448 lags = -6.26817163216166e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20217129491208+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 8.29468785234288e-9   nfactor = {1.98092133839856+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -4.50377981622488e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.409355e-05 letab = -3.95779542849e-11 petab = 6.16297582203915e-33   dsub = -0.0709802236591202 ldsub = 2.1852786982936e-7   voffl = 0.0   minv = 0.0   pclm = 0.61256302867136 lpclm = 7.68784699488308e-9   pdiblc1 = -0.22851602786032 lpdiblc1 = 2.15866014935975e-7   pdiblc2 = -0.012642675390946 lpdiblc2 = 7.41268117976658e-9   pdiblcb = 0.2251104 lpdiblcb = -1.407216152352e-07 wpdiblcb = -2.64697796016969e-23   drout = 1.71071422536632 ldrout = -3.99874830331655e-7   pscbe1 = 800088964.26928 lpscbe1 = -0.0500546785392544   pscbe2 = 9.4515592034632e-09 lpscbe2 = -7.56231627801261e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.70514182421279 lbeta0 = 1.8383773309196e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.26475020007599e-10 lagidl = -1.95859897305136e-16   bgidl = 653150899.0464 lbgidl = 195.150484462331   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.503945507280001 lkt1 = -2.54002515499539e-9   kt2 = -0.102203752992 lkt2 = 2.64528492319129e-8   at = 63054.141088 lat = 0.00109481416652982   ute = -0.30986055872 lute = 3.89517430971033e-8   ua1 = 7.4838232584e-10 lua1 = -1.08123453065966e-16   ub1 = 6.9220960552e-19 lub1 = -7.91629446505621e-26   uc1 = 5.401768370832e-11 luc1 = -1.67090453662817e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.70 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.09172011158686+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.14979819900128e-8   k1 = -1.32067307505343 lk1 = 5.94299434616013e-7   k2 = 0.661320056770371 lk2 = -2.14582026899029e-07 wk2 = -1.05879118406788e-22 pk2 = -2.52435489670724e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 13610.8058002857 lvsat = 0.0407792452282303   ua = 1.71355244464142e-09 lua = -1.02817043172251e-15   ub = -1.31803770378e-18 lub = 8.41818177747572e-25   uc = -5.466814300418e-13 luc = 1.88243636397102e-19 wuc = 1.92592994438724e-34 puc = 4.59177480789956e-41   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0118559007011428 lu0 = -2.3479741268039e-9   a0 = -0.140729426 la0 = 2.97893812465788e-7   keta = -0.138541690229726 lketa = 4.01965068889482e-08 wketa = -2.64697796016969e-23 pketa = 6.31088724176809e-30   a1 = 0.0   a2 = -0.0414961723505716 la2 = 1.76709072891218e-7   ags = -2.44893826583886 lags = 8.97502982946607e-7   b0 = 0.0   b1 = -7.30459064644572e-24 lb1 = 2.28369261052349e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0465650170048568+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.03537476600155e-8   nfactor = {5.77752696045714+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.2320009866314e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.45580506483057 leta0 = -3.019473638585e-7   etab = 0.109097785034743 letab = -3.41276531926919e-08 wetab = -2.52290086828673e-23 petab = -5.52202633654708e-30   dsub = 1.870698467732 ldsub = -3.88514672889777e-07 wdsub = -1.6940658945086e-21   voffl = 0.0   minv = 0.0   pclm = 0.689473970528859 lpclm = -1.63574360455608e-8   pdiblc1 = 1.535477391924 lpdiblc1 = -3.35625359838555e-7   pdiblc2 = 0.04140603300786 lpdiblc2 = -9.48499891661935e-9   pdiblcb = -0.744938571428571 lpdiblcb = 1.62552555094286e-7   drout = -1.538265090594 ldrout = 6.15879565051547e-7   pscbe1 = 799682270.466856 lpscbe1 = 0.0770932584628099   pscbe2 = 8.59036890806285e-09 lpscbe2 = 1.93617648793239e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 11.0290353605828 lbeta0 = -5.42699694331699e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 2228509545.27428 lbgidl = -297.366491977062   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.0752869374285723 lkt1 = -1.36554983116206e-7   kt2 = 0.337380461485714 lkt2 = -1.10977880413971e-7   at = 92247.8979428571 lat = -0.00803226358905895   ute = -0.0781973168571426 lute = -3.34749895124165e-8   ua1 = 1.27617545028571e-09 lua1 = -2.73131639906425e-16   ub1 = 4.39e-19   uc1 = -7.06743548285717e-13 luc1 = 3.99890122368949e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.71 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.26e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.0797208030717655+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.14051506229473e-07 wvth0 = -6.80183264231834e-07 pvth0 = 1.65038306866683e-13   k1 = 4.38070139821437 lk1 = -7.89070664828739e-07 wk1 = -5.40281734927562e-06 pk1 = 1.31092879599354e-12   k2 = -1.53238595079256 lk2 = 3.17694411364026e-07 wk2 = 2.18117756173318e-06 pk2 = -5.29236561223814e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 828523.074663173 lvsat = -0.156949437864123 wvsat = 0.0794741725403751 pvsat = -1.92834542768513e-8   ua = -6.60844309053298e-09 lua = 9.91061920941141e-16 wua = 3.919915287844e-15 pua = -9.51120405611895e-22   ub = 5.1528349803806e-18 lub = -7.28261428591789e-25 wub = -3.30212221451056e-24 pub = 8.01220329884413e-31   uc = 2.48548705198294e-12 luc = -5.47475659744416e-19 wuc = -2.09726024916604e-18 puc = 5.08875032337149e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00821545000223448 lu0 = 2.52209826516217e-09 wu0 = 8.8380914227875e-09 pu0 = -2.14445682664231e-15   a0 = -2.3714019079635 la0 = 8.39139722144445e-07 wa0 = 5.54234730716872e-06 pa0 = -1.3447840659168e-12   keta = 0.868810004974822 lketa = -2.04225293732093e-07 wketa = -5.95704321328443e-07 pketa = 1.44540505118491e-13   a1 = 0.0   a2 = 2.52175094444519 la2 = -4.45232081033874e-07 wa2 = -3.73156209201416e-06 pa2 = 9.05418762882131e-13   ags = 1.25   b0 = 0.0   b1 = 1.70440448417067e-23 lb1 = -3.62421160705082e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.870148199686177+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.59478828619415e-07 wvoff = 5.74922984701727e-07 pvoff = -1.39498163162058e-13   nfactor = {-12.8339372210939+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.28384745945179e-06 wnfactor = 7.22684153815738e-06 pnfactor = -1.75350637713543e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 3.52227140742454 leta0 = -8.03350624292817e-07 weta0 = -3.90426658603447e-06 peta0 = 9.47323435902232e-13   etab = 0.218998464849793 letab = -6.07937343416561e-08 wetab = -4.36768612044607e-07 petab = 1.05976662489279e-13   dsub = 0.494630368576166 ldsub = -5.46282614468046e-08 wdsub = -1.86483773502629e-07 pdsub = 4.52480498351311e-14   voffl = 0.0   minv = 0.0   pclm = -3.41874242342863 lpclm = 9.80451973351495e-07 wpclm = 4.82055278961276e-06 ppclm = -1.16964928776606e-12   pdiblc1 = -2.85585094980011 lpdiblc1 = 7.298777663407e-07 wpdiblc1 = 3.63716160230719e-06 ppdiblc1 = -8.82513616860613e-13   pdiblc2 = -0.0558310351752088 lpdiblc2 = 1.41084088331841e-08 wpdiblc2 = 6.5859884998796e-08 ppdiblc2 = -1.59801107763379e-14   pdiblcb = 4.28307778464816 lpdiblcb = -1.05743527751146e-06 wpdiblcb = -4.50343559687385e-06 ppdiblcb = 1.09270460635428e-12   drout = 1.0   pscbe1 = 800000000.0   pscbe2 = 1.5828270404401e-08 lpscbe2 = -1.56257229447526e-15 wpscbe2 = -5.85177821868213e-15 ppscbe2 = 1.41986376342459e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -2.40008019514829 lbeta0 = 2.71571404587977e-06 wbeta0 = 2.03697256529492e-05 pbeta0 = -4.9424694929803e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.10020582196878e-08 lagidl = -2.64525360230862e-15 wagidl = -1.53937456985719e-14 pagidl = 3.7351076688101e-21   bgidl = 1023886902.30666 lbgidl = -5.07926313268581   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.130016938666664 lkt1 = -1.23275405075797e-7   kt2 = -0.12   at = -631791.338530377 lat = 0.167647168670334 wat = 0.884683951267534 pat = -2.14657944567652e-7   ute = -0.242597991333333 lute = 6.4148613411373e-9   ua1 = -1.97352441537341e-09 lua1 = 5.15369036097374e-16 wua1 = 2.23624901166777e-15 pua1 = -5.42598987693046e-22   ub1 = 9.35793247333334e-19 lub1 = -1.20540919946466e-25   uc1 = -1.12695701272335e-13 luc1 = 2.55751540865296e-19 wuc1 = -4.48554602181233e-17 puc1 = 1.0883639156405e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.72 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.003036+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.010197753   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.38874612e-9   ub = 1.066826e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0048880282   a0 = 1.279916   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21647917   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17570541+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4613328+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.73 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.003036+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.49177002   k2 = 0.010197753   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55237.817   ua = -1.38874612e-9   ub = 1.066826e-18   uc = -3.8916596e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0048880282   a0 = 1.279916   keta = 0.0066402373   a1 = 0.0   a2 = 0.8   ags = 0.21647917   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17570541+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.4613328+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00056783834   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799985290.0   pscbe2 = 1.0771971e-8   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.4670794e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.54561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.74 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.981642148292+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.72490881747283e-7   k1 = 0.534439388927654 lk1 = -3.44027675352131e-7   k2 = 0.005689110475084 lk2 = 3.63515525498037e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 67925.4832099965 lvsat = -0.102296059716033   ua = -2.02129883628681e-09 lua = 5.10004356733725e-15   ub = 1.52617076555832e-18 lub = -3.7035305618916e-24   uc = -2.30174367955125e-11 luc = -1.28189165170151e-16   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0026427586981379 lu0 = 1.81027952059544e-8   a0 = 1.341190737635 la0 = -4.94036028095985e-7   keta = 0.0101116040437775 lketa = -2.79883734203168e-08 wketa = -6.61744490042422e-24   a1 = 0.0   a2 = 0.8   ags = 0.170330354757245 lags = 3.72081191431215e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.174175329119845+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.23364882474125e-8   nfactor = {0.315488909136601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.23852449654312e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.0350910319060362 lpclm = 2.96957167307167e-07 wpclm = -3.30872245021211e-24 ppclm = -2.52435489670724e-29   pdiblc1 = 0.39   pdiblc2 = 9.04296639703799e-05 lpdiblc2 = 3.8491733328861e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799970369.961945 lpscbe1 = 0.12029486578831   pscbe2 = 1.20609351273826e-08 lpscbe2 = -1.03924511540718e-14   pvag = 0.0   delta = 0.01   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.35768627006325e-10 lagidl = 8.81997206366977e-17   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.631260565635 lkt1 = 6.90569505210245e-7   kt2 = -0.078629106849 lkt2 = 2.10798531994808e-7   at = -35977.38207575 lat = 0.370698987864461 pat = 5.29395592033938e-23   ute = -2.46762697525 lute = 9.74069045947571e-6   ua1 = -2.465769591175e-09 lua1 = 1.7816169145152e-14 wua1 = 3.94430452610506e-31 pua1 = -6.01853107621011e-36   ub1 = 2.02782333948e-18 lub1 = -1.23639210452584e-23 pub1 = -2.80259692864963e-45   uc1 = 9.77712911684499e-11 luc1 = -7.22220402810009e-16 wuc1 = 1.23259516440783e-32 puc1 = -1.41059322098675e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.75 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0166179869188+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.03967106601799e-8   k1 = 0.437921473358791 lk1 = 4.80896761187344e-8   k2 = 0.01471198164958 lk2 = -3.05106752808383e-10   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 31719.18570813 lvsat = 0.0447970203543542   ua = -5.02669836569194e-10 lua = -1.06959631481753e-15   ub = 4.6494729061422e-19 lub = 6.07836253908345e-25   uc = -6.4407623172087e-11 luc = 3.99641788304033e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0081896092382 lu0 = -4.43205057842235e-9   a0 = 1.3104492260441 la0 = -3.69144394929349e-7   keta = 0.0115107076952954 lketa = -3.36724250809121e-08 pketa = 1.26217744835362e-29   a1 = 0.0   a2 = 0.8   ags = 0.14144178625091 lags = 4.89444987610655e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.17061466580209+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.68021743473283e-8   nfactor = {3.6130470793536+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.15826063299095e-06 wnfactor = 3.3881317890172e-21   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.1619898605 leta0 = -3.33095122881999e-7   etab = -0.141676668963335 letab = 2.91196359043864e-7   dsub = 0.8693957 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = -0.286123216206924 lpclm = 1.31681005847096e-06 wpclm = 1.05879118406788e-22 ppclm = -4.03896783473158e-28   pdiblc1 = 0.39   pdiblc2 = 0.0018865445760297 lpdiblc2 = -3.44779136121275e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 799999959.37362 lpscbe1 = 8.37975130707491e-5   pscbe2 = 9.63772154963349e-09 lpscbe2 = -5.47811590992355e-16   pvag = 0.0   delta = 0.01   alpha0 = -3.144478223853e-12 lalpha0 = 1.27748767223977e-17   alpha1 = 3.0154328869995e-15 lalpha1 = -1.22506122331739e-20   beta0 = 57.845613 lbeta0 = -0.000113126645507094   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.37277016954701e-11 lagidl = 3.80875921359739e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.45128651889 lkt1 = -4.05998961097684e-8   kt2 = -0.007366609947 lkt2 = -7.87151958941399e-8   at = 104574.830071 lat = -0.200313770186987   ute = 0.78088974095 lute = -3.45685699539363e-06 wute = -1.05879118406788e-22 pute = -4.03896783473158e-28   ua1 = 4.05743146829e-09 lua1 = -8.68523536067075e-15   ub1 = -2.83288002861e-18 lub1 = 7.38335716467207e-24   uc1 = -2.26309101254e-10 luc1 = 5.94400914500348e-16 puc1 = 1.88079096131566e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.76 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0393498757844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.64909471257836e-8   k1 = 0.469339308574519 lk1 = -1.67139446749709e-8   k2 = 0.021958720811088 lk2 = -1.52525063234229e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 79606.936194042 lvsat = -0.0539780735324065   ua = -1.32936764173355e-09 lua = 6.35581992631081e-16   ub = 9.34438395790239e-19 lub = -3.60553940289709e-25   uc = -4.11564853467139e-11 luc = -7.99450159144852e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0045993584211 lu0 = 2.97333718645915e-9   a0 = 1.5849937892658 la0 = -9.3543044372383e-7   keta = 0.0302810020398646 lketa = -7.23887474672056e-08 pketa = 2.52435489670724e-29   a1 = 0.0   a2 = 0.8   ags = -0.372591207902342 lags = 1.54970897460493e-06 pags = -4.03896783473158e-28   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1677958864496+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.26162957533895e-8   nfactor = {1.2213286935428+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.74988594881063e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.083979721 leta0 = 1.74251082763998e-07 weta0 = 6.61744490042422e-24 peta0 = -2.68212707775144e-29   etab = 0.00640714392666938 letab = -1.42469406079481e-08 petab = -5.52202633654708e-30   dsub = -0.0587914000000005 ldsub = 6.575512557132e-7   voffl = 0.0   minv = 0.0   pclm = 0.33200266945972 lpclm = 4.18401179112811e-8   pdiblc1 = 0.39824678284746 lpdiblc1 = -1.70101276789189e-8   pdiblc2 = 0.000215   pdiblcb = -0.4375276 lpdiblcb = 4.383675038088e-7   drout = 0.186745427113599 ldrout = 7.69889065709258e-7   pscbe1 = 800000000.0   pscbe2 = 1.039468368145e-08 lpscbe2 = -2.10915044863806e-15   pvag = 0.0   delta = 0.01   alpha0 = -9.99748435522941e-11 lalpha0 = 2.12500867802723e-16 walpha0 = 2.46519032881566e-32 palpha0 = 5.87747175411144e-38   alpha1 = -1.06269830865774e-10 lalpha1 = 2.19190160531544e-16 walpha1 = -2.6638018543306e-32 palpha1 = 1.40278720381332e-38   beta0 = -3.27065467911561 lbeta0 = 1.29340906260216e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.0605930052948e-10 lagidl = -3.25230242996046e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.42540755738626 lkt1 = -9.39788255079199e-8   kt2 = -0.0260334075704199 lkt2 = -4.02123497777639e-8   at = -9001.35875991802 lat = 0.0339527927908397   ute = -0.577978479603001 lute = -6.54003766688627e-7   ua1 = -6.069851608966e-11 lua1 = -1.91023965949856e-16   ub1 = 1.03017017304036e-18 lub1 = -5.84716977159622e-25   uc1 = 7.71992542605119e-11 luc1 = -3.1626952901394e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.77 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.05137782399656+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.9272301958057e-8   k1 = 0.391153407181879 lk1 = 6.63693652091016e-8   k2 = 0.0238942373178024 lk2 = -1.73092597130849e-08 pk2 = 6.31088724176809e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -23746.9038300841 lvsat = 0.0558496443231508   ua = -2.80252503543959e-10 lua = -4.79247619584434e-16   ub = 2.12775299295278e-19 lub = 4.06312689243502e-25   uc = -7.89302775186919e-11 luc = 3.21453653745978e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00867088346895599 lu0 = -1.35322004734446e-9   a0 = 0.220162530228 la0 = 5.14891115717578e-7   keta = -0.042886499465348 lketa = 5.36181999729047e-9   a1 = 0.0   a2 = 0.8   ags = 0.830448601759198 lags = 2.71313157345808e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.21093603152804+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.32260617324734e-8   nfactor = {2.00663010659672+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.95025280837248e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.38136316 leta0 = 4.9026202561608e-07 weta0 = 1.05879118406788e-22 peta0 = -1.0097419586829e-28   etab = -0.014869899025 letab = 8.36285376012795e-9   dsub = 0.832971162499519 ldsub = -2.90069530176164e-7   voffl = 0.0   minv = 0.0   pclm = 0.0845993725202803 lpclm = 3.04740262564414e-7   pdiblc1 = 0.637775646199679 lpdiblc1 = -2.71542599973796e-7   pdiblc2 = -0.000141928826311 lpdiblc2 = 3.79286134133468e-10   pdiblcb = -0.025   drout = 0.8113877057728 ldrout = 1.06120443999403e-7   pscbe1 = 800000000.0   pscbe2 = 7.38890444982519e-09 lpscbe2 = 1.08490478249725e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.7537747206644 lbeta0 = 1.56475017498226e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.132375100038e-10 lagidl = 3.32858081155418e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.519908287987479 lkt1 = 6.44124185669976e-9   kt2 = -0.0736511439751598 lkt2 = 1.03880663998961e-8   at = -24367.726158164 lat = 0.0502816787101771   ute = -2.265596160714 lute = 1.1393229107318e-6   ua1 = -1.13693879534068e-09 lua1 = 9.5262985191289e-16 pua1 = -3.76158192263132e-37   ub1 = 3.99361023599279e-19 lub1 = 8.56047957841481e-26   uc1 = 7.34491041749761e-11 luc1 = -2.76419009148001e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.78 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.00983041569376+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.89615124538495e-9   k1 = 0.420161160566559 lk1 = 5.00485008602523e-8   k2 = 0.0158511726935312 lk2 = -1.27839259190142e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -10183.06594408 lvsat = 0.0482181137026452   ua = -5.77918020554799e-10 lua = -3.11769688424489e-16   ub = 3.85114607900799e-19 lub = 3.0934804532831e-25   uc = -4.91245534217428e-11 luc = 1.53755323801385e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.008666870117048 lu0 = -1.35096198305365e-9   a0 = 1.53946590088 la0 = -2.27399094139322e-7   keta = -0.0626034569112048 lketa = 1.64553295007124e-8   a1 = 0.0   a2 = 1.14549842976048 la2 = -1.94390545523577e-7   ags = 2.42673310540448 lags = -6.26817163216166e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20217129491208+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 8.29468785234288e-9   nfactor = {1.98092133839856+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -4.5037798162248e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.409355e-05 letab = -3.95779542849e-11 wetab = -1.29246970711411e-26 petab = 3.08148791101958e-33   dsub = -0.0709802236591193 ldsub = 2.1852786982936e-7   voffl = 0.0   minv = 0.0   pclm = 0.61256302867136 lpclm = 7.68784699488393e-9   pdiblc1 = -0.228516027860321 lpdiblc1 = 2.15866014935975e-07 ppdiblc1 = -1.0097419586829e-28   pdiblc2 = -0.012642675390946 lpdiblc2 = 7.41268117976657e-09 ppdiblc2 = 5.91645678915759e-31   pdiblcb = 0.2251104 lpdiblcb = -1.407216152352e-07 wpdiblcb = 5.29395592033938e-23   drout = 1.71071422536632 ldrout = -3.99874830331655e-7   pscbe1 = 800088964.269281 lpscbe1 = -0.0500546785392544   pscbe2 = 9.45155920346318e-09 lpscbe2 = -7.56231627801198e-17   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.7051418242128 lbeta0 = 1.83837733091957e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 7.264750200076e-10 lagidl = -1.95859897305136e-16   bgidl = 653150899.0464 lbgidl = 195.150484462331   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.503945507279999 lkt1 = -2.54002515499539e-9   kt2 = -0.102203752992 lkt2 = 2.64528492319129e-8   at = 63054.1410879999 lat = 0.00109481416652984   ute = -0.30986055872 lute = 3.89517430971034e-8   ua1 = 7.4838232584e-10 lua1 = -1.08123453065966e-16   ub1 = 6.9220960552e-19 lub1 = -7.91629446505617e-26   uc1 = 5.401768370832e-11 luc1 = -1.67090453662818e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.79 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.09172011158686+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.14979819900111e-8   k1 = -1.32067307505343 lk1 = 5.94299434616013e-7   k2 = 0.661320056770372 lk2 = -2.14582026899029e-07 wk2 = -1.05879118406788e-22 pk2 = -2.52435489670724e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 13610.8058002861 lvsat = 0.0407792452282304   ua = 1.71355244464142e-09 lua = -1.02817043172251e-15   ub = -1.31803770378e-18 lub = 8.41818177747569e-25   uc = -5.466814300418e-13 luc = 1.88243636397102e-19 puc = 4.59177480789956e-41   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0118559007011429 lu0 = -2.3479741268039e-9   a0 = -0.140729426 la0 = 2.97893812465788e-7   keta = -0.138541690229726 lketa = 4.01965068889482e-08 wketa = -5.29395592033938e-23   a1 = 0.0   a2 = -0.0414961723505698 la2 = 1.76709072891218e-7   ags = -2.44893826583886 lags = 8.9750298294661e-7   b0 = 0.0   b1 = -7.30459064644571e-24 lb1 = 2.28369261052349e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0465650170048573+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.03537476600156e-8   nfactor = {5.77752696045714+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.2320009866314e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.45580506483057 leta0 = -3.019473638585e-7   etab = 0.109097785034743 letab = -3.41276531926919e-08 wetab = -3.66027421054715e-23 petab = -4.33873497871556e-30   dsub = 1.870698467732 ldsub = -3.88514672889777e-07 wdsub = 1.6940658945086e-21   voffl = 0.0   minv = 0.0   pclm = 0.689473970528857 lpclm = -1.63574360455608e-8   pdiblc1 = 1.535477391924 lpdiblc1 = -3.35625359838555e-7   pdiblc2 = 0.04140603300786 lpdiblc2 = -9.48499891661934e-9   pdiblcb = -0.744938571428571 lpdiblcb = 1.62552555094286e-7   drout = -1.538265090594 ldrout = 6.15879565051547e-7   pscbe1 = 799682270.466858 lpscbe1 = 0.0770932584628099   pscbe2 = 8.59036890806285e-09 lpscbe2 = 1.93617648793245e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 11.0290353605829 lbeta0 = -5.42699694331699e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.0e-10   bgidl = 2228509545.27428 lbgidl = -297.366491977062   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.0752869374285705 lkt1 = -1.36554983116207e-7   kt2 = 0.337380461485714 lkt2 = -1.10977880413971e-07 wkt2 = -5.29395592033938e-23 pkt2 = -1.26217744835362e-29   at = 92247.8979428571 lat = -0.00803226358905895   ute = -0.0781973168571435 lute = -3.34749895124164e-8   ua1 = 1.27617545028571e-09 lua1 = -2.73131639906425e-16   ub1 = 4.39e-19   uc1 = -7.06743548285713e-13 luc1 = 3.99890122368949e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.80 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-2.05298032517951+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.64736237695708e-07 wvth0 = 1.13727202718124e-06 pvth0 = -2.75945410131203e-13   k1 = -6.76709541112815 lk1 = 1.91580845739651e-06 wk1 = 4.86477394915419e-06 pk1 = -1.18037902147488e-12   k2 = 2.69381299145171 lk2 = -7.07742047584239e-07 wk2 = -1.71133000966916e-06 pk2 = 4.15233690886105e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 951996.675552068 lvsat = -0.186908825436603 wvsat = -0.0342502244642562 pvsat = 8.31040596355793e-9   ua = 1.32064560017303e-08 lua = -3.81678556500743e-15 wua = -1.43304429648722e-14 pua = 3.47711002011065e-21   ub = -1.40572506736061e-17 lub = 3.93283533432023e-24 wub = 1.43911773384258e-23 pub = -3.49184648704095e-30   uc = -2.40934195906179e-12 luc = 6.40195861837454e-19 wuc = 2.41108383179042e-18 puc = -5.85020558777965e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0368024340507847 lu0 = -8.4009510856943e-09 wu0 = -3.26252795447502e-08 pu0 = 7.91613257817911e-15   a0 = 14.478638439623 la0 = -3.24932036771325e-06 wa0 = -9.97725092466114e-06 pa0 = 2.42086020985793e-12   keta = 3.49264746559229 lketa = -8.40867967501394e-07 wketa = -3.01236934849797e-06 pketa = 7.3091527398085e-13   a1 = 0.0   a2 = -1.52970521251935 la2 = 5.37805137979686e-7   ags = -21.3748093653398 lags = 5.48963849478733e-06 wags = 2.08384041924332e-05 pags = -5.05618871644361e-12   b0 = 0.0   b1 = 1.70440448417067e-23 lb1 = -3.62421160705082e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.667379380948574+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.10279407978561e-07 wvoff = 3.88164345800247e-07 pvoff = -9.41834205362804e-14   nfactor = {-32.0405360913802+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 7.94409819614031e-06 wnfactor = 2.49169296161634e-05 pnfactor = -6.04579396820665e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.28176546236366 leta0 = -2.59718742795135e-07 weta0 = -1.84066606128252e-06 peta0 = 4.46615531777468e-13   etab = -1.65477112576423 letab = 3.9385397158575e-07 wetab = 1.28905225398763e-06 petab = -3.12773060803052e-13   dsub = 0.0801490693944764 ldsub = 4.5940652024043e-08 wdsub = 1.95270994154533e-07 pdsub = -4.73801634796676e-14   voffl = 0.0   minv = 0.0   pclm = -3.86271696503177 lpclm = 1.088177068177e-06 wpclm = 5.22947207815491e-06 ppclm = -1.26886864609935e-12   pdiblc1 = 1.09311208610333 lpdiblc1 = -2.2829072676484e-7   pdiblc2 = 0.01567479267806 lpdiblc2 = -3.24162222547732e-9   pdiblcb = -0.60642195474906 lpdiblcb = 1.28943160256403e-7   drout = 1.0   pscbe1 = -243568471.767365 lpscbe1 = 253.209366852688 wpscbe1 = 961.170601087244 ppscbe1 = -0.000233216512306606   pscbe2 = -9.89944972601599e-09 lpscbe2 = 4.67995026252885e-15 wpscbe2 = 1.78445377312213e-14 ppscbe2 = -4.32976294602808e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 20.0381566215414 lbeta0 = -2.72865485884814e-06 wbeta0 = -2.9683734881561e-07 pbeta0 = 7.20240206419156e-14   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.92610521695205e-08 lagidl = 7.12410697630811e-15 wagidl = 2.16902780731473e-14 pagidl = -5.26288569111233e-21   bgidl = 1023886902.30666 lbgidl = -5.07926313268763   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.130016938666664 lkt1 = -1.23275405075797e-7   kt2 = -0.12   at = 328733.544333334 lat = -0.0654126678579513   ute = -0.242597991333332 lute = 6.41486134113751e-9   ua1 = 4.54430581333332e-10 lua1 = -7.37451083935573e-17   ub1 = 9.35793247333331e-19 lub1 = -1.20540919946465e-25   uc1 = -4.88134612233334e-11 luc1 = 1.20724078856072e-17 wuc1 = -6.16297582203915e-33 puc1 = 1.46936793852786e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.81 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.905187715630101+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -7.44666736030938e-8   k1 = 0.52852970130877 wk1 = -2.79756687345252e-8   k2 = -0.00276816367190749 wk2 = 9.86760974900517e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 141489.070159167 wvsat = -0.0656408434570094   ua = -2.75554094157253e-09 wua = 1.04018853795817e-15   ub = 2.07757424036045e-18 wub = -7.69222064490046e-25   uc = 4.2695284193716e-11 wuc = -6.21100848487621e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.000160468239056095 wu0 = 3.84211883667142e-9   a0 = 1.3612227966662 wa0 = -6.18779034097977e-8   keta = 0.0044876067427465 wketa = 1.63824269507943e-9   a1 = 0.0   a2 = 0.8   ags = 0.16462801455343 wags = 3.94609174135996e-8   b0 = 9.1668685058e-08 wb0 = -6.97637377476475e-14   b1 = -5.3498178981e-09 wb1 = 4.0714371827694e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.13423864073745+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -3.15579613064634e-8   nfactor = {1.6634485330711+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.53818602151042e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = -0.00018967155319159 wpdiblc2 = 5.76496995636293e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 827723160.26378 wpscbe1 = -21.1096898088613   pscbe2 = 1.42901336691986e-08 wpscbe2 = -2.67747025772477e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.805211e-10 walpha0 = 2.1348839509042e-16   alpha1 = -2.805211e-10 walpha1 = 2.1348839509042e-16   beta0 = 105.740697 wbeta0 = -5.76418666744134e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.73272686720386e-09 wagidl = 2.191371400431e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60171422 wkt1 = 4.26976790180839e-8   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.82 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.905187715630101+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -7.44666736030938e-8   k1 = 0.52852970130877 wk1 = -2.7975668734525e-8   k2 = -0.00276816367190749 wk2 = 9.86760974900515e-9   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 141489.070159167 wvsat = -0.0656408434570094   ua = -2.75554094157253e-09 wua = 1.04018853795817e-15   ub = 2.07757424036045e-18 wub = -7.69222064490046e-25   uc = 4.2695284193716e-11 wuc = -6.2110084848762e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.000160468239056095 wu0 = 3.84211883667142e-9   a0 = 1.3612227966662 wa0 = -6.18779034097964e-8   keta = 0.00448760674274651 wketa = 1.63824269507943e-9   a1 = 0.0   a2 = 0.8   ags = 0.16462801455343 wags = 3.94609174135996e-8   b0 = 9.1668685058e-08 wb0 = -6.97637377476475e-14   b1 = -5.3498178981e-09 wb1 = 4.0714371827694e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.13423864073745+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -3.15579613064634e-8   nfactor = {1.6634485330711+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.53818602151043e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = -0.00018967155319159 wpdiblc2 = 5.76496995636292e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 827723160.263781 wpscbe1 = -21.1096898088617   pscbe2 = 1.42901336691986e-08 wpscbe2 = -2.67747025772477e-15   pvag = 0.0   delta = 0.01   alpha0 = -2.805211e-10 walpha0 = 2.1348839509042e-16   alpha1 = -2.805211e-10 walpha1 = 2.1348839509042e-16   beta0 = 105.740697 wbeta0 = -5.76418666744134e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.73272686720386e-09 wagidl = 2.191371400431e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60171422 wkt1 = 4.26976790180839e-8   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.83 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.777253722443274+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.03148547495986e-06 wvth0 = -1.55548217262453e-07 pvth0 = 6.53731135006601e-13   k1 = 0.644515798364248 lk1 = -9.35153913591186e-07 wk1 = -8.37727928057256e-08 pk1 = 4.49872012827175e-13   k2 = -9.94156963803616e-05 lk2 = -2.15171488399081e-08 wk2 = 4.40531269228882e-09 pk2 = 4.40405238167694e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 279416.425183049 lvsat = -1.11205833385504 wvsat = -0.160953531759244 pvsat = 7.68471702587753e-7   ua = -5.02429572306754e-09 lua = 1.82921485139633e-14 wua = 2.28540735730875e-15 pua = -1.00397485712112e-20   ub = 3.56022951745317e-18 lub = -1.19541127779883e-23 wub = -1.54800454747131e-24 pub = 6.27904124101909e-30   uc = 8.98817299030025e-11 luc = -3.80447230260631e-16 wuc = -8.59210302024046e-17 puc = 1.91979032824202e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00761412118911264 lu0 = 6.0096105513938e-08 wu0 = 7.8059184345289e-09 pu0 = -3.19586812620705e-14   a0 = 1.58592244942458 la0 = -1.81167195891653e-06 wa0 = -1.86251160350108e-07 pa0 = 1.00277654759072e-12   keta = 0.0269043821605375 lketa = -1.80738345320948e-07 wketa = -1.27800128020909e-08 pketa = 1.16249174665194e-13   a1 = 0.0   a2 = 0.8   ags = -0.0136050136461545 lags = 1.43702838601704e-06 wags = 1.39982577427534e-07 pags = -8.10469755851426e-13   b0 = 1.00506714861532e-07 lb0 = -7.12578349390918e-14 wb0 = -7.64898513929932e-14 pb0 = 5.42302194692833e-20   b1 = -1.03137591635746e-08 lb1 = 4.00224614767834e-14 wb1 = 7.84920596411695e-15 pb1 = -3.04587821317065e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0992837693475173+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.81828474353586e-07 wvoff = -5.69956374105639e-08 pvoff = 2.05094773988612e-13   nfactor = {-1.28052671099136+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.37362066738373e-05 wnfactor = 1.21463523877654e-06 pnfactor = -1.10333479391087e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.995801739932209 lpclm = -8.0147580688412e-06 wpclm = -7.84552903043876e-07 ppclm = 6.32556604909187e-12   pdiblc1 = 0.39   pdiblc2 = -0.00316840503606394 lpdiblc2 = 2.4016449770879e-08 wpdiblc2 = 2.48011072955046e-09 ppdiblc2 = -1.53481484283783e-14   pdiblcb = -0.225   drout = 0.56   pscbe1 = 855880528.651685 lpscbe1 = -227.022668344322 wpscbe1 = -42.5499901715884 ppscbe1 = 0.000172865380435936   pscbe2 = 1.93701874907277e-08 lpscbe2 = -4.09586349835054e-14 wpscbe2 = -5.56264949895532e-15 ppscbe2 = 2.32621557871566e-20   pvag = 0.0   delta = 0.01   alpha0 = -5.04798893201368e-10 lalpha0 = 1.80827065802149e-15 walpha0 = 3.84173260239534e-16 palpha0 = -1.37617027977612e-21   alpha1 = -5.65434924367384e-10 lalpha1 = 2.2971570270698e-15 walpha1 = 4.30319838797387e-16 palpha1 = -1.74823343762666e-21   beta0 = 164.620583219651 lbeta0 = -0.000474727208070234 wbeta0 = -0.000102451944818766 pbeta0 = 3.61287438829628e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -5.83195600078963e-09 lagidl = 2.49879625831557e-14 wagidl = 4.54169027973201e-15 pagidl = -1.89497703083698e-20   bgidl = 1916374054.79262 lbgidl = -7388.39227638506 wbgidl = -697.399326682296 pbgidl = 0.0056228783124831   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.549665888019039 lkt1 = -4.1964685926632e-07 wkt1 = -6.20969929611426e-08 pkt1 = 8.44921504497247e-13   kt2 = -0.169190893900297 lkt2 = 9.409654376225e-07 wkt2 = 6.89213416534503e-08 pkt2 = -5.55687828226091e-13   at = -14516.2040004778 lat = 0.197665277990005 wat = -0.0163328621769969 pat = 1.31685955237018e-7   ute = -3.30484652965617 lute = 1.6490888653174e-05 wute = 6.37159411568295e-07 pute = -5.13718568376818e-12   ua1 = -6.86737625241902e-09 lua1 = 5.33047302731512e-14 wua1 = 3.3498084170078e-15 pua1 = -2.7008292635687e-20   ub1 = 6.12723673509394e-18 lub1 = -4.54160072664444e-23 wub1 = -3.11982658930751e-24 pub1 = 2.51540324123611e-29   uc1 = 1.9920328789939e-10 luc1 = -1.54002987406876e-15 wuc1 = -7.71940299425075e-17 puc1 = 6.22387519187599e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.84 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.09565134754287+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.62048815879536e-07 wvth0 = 6.01477226427385e-08 pvth0 = -2.22563386897944e-13   k1 = 0.33180900427363 lk1 = 3.35260590939536e-07 wk1 = 8.07560669200021e-08 pk1 = -2.18549184791236e-13   k2 = -0.0252653029596089 lk2 = 8.07227410594e-08 wk2 = 3.04244006290032e-08 pk2 = -6.16656115602682e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -104730.891711536 lvsat = 0.448593153358942 wvsat = 0.103844267109633 pvsat = -3.07305897413304e-7   ua = 1.40909812711933e-09 lua = -7.84440181077216e-15 wua = -1.45493609697504e-15 pua = 5.15591287921341e-21   ub = -5.32183992536304e-19 lub = 4.67188185940833e-24 wub = 7.58858985417698e-25 pub = -3.09291020851004e-30   uc = -2.30768246133936e-11 luc = 7.84624857427521e-17 wuc = -3.14544818628649e-17 puc = -2.92988361888492e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0153062323647307 lu0 = -3.30209938073412e-08 wu0 = -5.41605052078584e-09 pu0 = 2.17573922506115e-14   a0 = 1.23647116492131 la0 = -3.91977891344723e-07 wa0 = 5.63004263886232e-08 pa0 = 1.73772543456451e-14   keta = -0.0321726784224514 lketa = 5.92703659318054e-08 wketa = 3.32449002744995e-08 pketa = -7.07333861464588e-14   a1 = 0.0   a2 = 0.8   ags = 0.855777420650232 lags = -2.09495772808796e-06 wags = -5.43639562741656e-07 pags = 1.96683952844125e-12   b0 = 1.67953292476843e-07 lb0 = -3.45268864129001e-13 wb0 = -1.2781954320382e-13 pb0 = 2.62764175948236e-19   b1 = -7.12704707637278e-10 lb1 = 1.01685280402319e-15 wb1 = 5.42398358650631e-16 pb1 = -7.73867895049974e-22   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.175226034731536+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.66974588016138e-08 wvoff = 3.50944635507707e-09 pvoff = -4.07154785108642e-14   nfactor = {9.87766277625092+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.15954779482338e-05 wnfactor = -4.76763691212127e-06 pnfactor = 1.32704582274705e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.1619898605 leta0 = -3.33095122881999e-7   etab = -0.141676664652664 letab = 2.91196341531171e-07 wetab = -3.28060212103357e-15 petab = 1.33278987482499e-20   dsub = 0.8693957 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = -2.49724551435336 lpclm = 6.17622844221503e-06 wpclm = 1.68275737825042e-06 ppclm = -3.69822245748503e-12   pdiblc1 = 0.39   pdiblc2 = 0.00556424430506413 lpdiblc2 = -1.14611432830629e-08 wpdiblc2 = -2.79888469272377e-09 ppdiblc2 = 6.09849897597909e-15   pdiblcb = 0.353613480661799 lpdiblcb = -2.35069711384889e-06 wpdiblcb = -4.40349276272513e-07 ppdiblcb = 1.78897970305721e-12   drout = 0.56   pscbe1 = 799999845.408051 lpscbe1 = 0.000318867227178998 wpscbe1 = 8.67326066327223e-05 ppscbe1 = -1.78897970222469e-10   pscbe2 = 9.65356460819317e-09 lpscbe2 = -1.48351362925122e-15 wpscbe2 = -1.20572361409873e-17 ppscbe2 = 7.12108737741027e-22   pvag = 0.0   delta = 0.01   alpha0 = -1.22490039814423e-10 lalpha0 = 2.55088182515259e-16 walpha0 = 9.08270087531227e-17 palpha0 = -1.84410651329872e-22   alpha1 = 9.81242463029571e-15 lalpha1 = -4.02475214397213e-20 walpha1 = -5.17279754969999e-21 palpha1 = 2.13068293757511e-26   beta0 = 93.9393574500413 lbeta0 = -0.000187574974372038 wbeta0 = -2.74688626824972e-05 pbeta0 = 5.66583199857007e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.9090307046073e-10 lagidl = -1.51205254835072e-15 wagidl = -4.77306922430925e-16 pagidl = 1.44059844703108e-21   bgidl = -832748109.585239 lbgidl = 3780.29589525868 wbgidl = 1394.79865336459 pbgidl = -0.00287696470477864   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.897859537891015 lkt1 = 9.94937894062268e-07 wkt1 = 3.39860912841174e-07 pkt1 = -7.88087958015665e-13   kt2 = 0.139122697421969 lkt2 = -3.11601074399807e-07 wkt2 = -1.11484544756556e-07 pkt2 = 1.77235981326886e-13   at = 155601.591821289 lat = -0.493461743791746 wat = -0.0388335190213157 pat = 2.23097978757708e-7   ute = 2.25173247148997 lute = -6.08348034688437e-06 wute = -1.11937338750415e-06 pute = 1.99897121398989e-12   ua1 = 1.32785125592757e-08 lua1 = -2.85407231570148e-14 wua1 = -7.01763183986218e-15 pua1 = 1.51108641146028e-20   ub1 = -1.16984235764688e-17 lub1 = 2.70031976904024e-23 wub1 = 6.74705276585829e-24 pub1 = -1.4931526597351e-29   uc1 = -4.74687560157723e-10 luc1 = 1.19774469310029e-15 wuc1 = 1.89026488796699e-16 puc1 = -4.59170076622014e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.85 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.904696002702602+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.31822934691114e-07 wvth0 = -1.02477279808692e-07 pvth0 = 1.12873122908472e-13   k1 = 0.631103332077813 lk1 = -2.8207526277383e-07 wk1 = -1.23109248327798e-07 pk1 = 2.01951161320856e-13   k2 = 0.0761814188385838 lk2 = -1.28525122296981e-07 wk2 = -4.12657613967811e-08 pk2 = 8.62052408602714e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 373263.725461541 lvsat = -0.5373367078177 wvsat = -0.223485208949074 pvsat = 3.67856318425475e-7   ua = -6.8857440504819e-09 lua = 9.26485486875089e-15 wua = 4.22863692614194e-15 pua = -6.56724081404254e-21   ub = 4.69092187832859e-18 lub = -6.10149478786069e-24 wub = -2.85884245381465e-24 pub = 4.36909825270528e-30   uc = 1.5304612735833e-10 luc = -2.84815407666299e-16 wuc = -1.47796383618794e-16 puc = 2.10672391365197e-22   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.0193982819600957 lu0 = 3.85618562105901e-08 wu0 = 1.8263217030514e-08 pu0 = -2.70843648128664e-14   a0 = 2.94980472092034 la0 = -3.92596479062345e-06 wa0 = -1.03867871401042e-06 pa0 = 2.27592283854005e-12   keta = 0.14769121136057 lketa = -3.11723727962466e-07 wketa = -8.93541240038898e-08 pketa = 1.8214402009307e-13   a1 = 0.0   a2 = -0.392369522647201 la2 = 2.45942668745398e-06 wa2 = 9.07443524728375e-07 pa2 = -1.87172749695869e-12   ags = -3.37354922400818 lags = 6.62861212359697e-06 wags = 2.28385569068482e-06 pags = -3.86525962609583e-12   b0 = 1.87564087558092e-07 lb0 = -3.85718835273799e-13 wb0 = -1.42744185836203e-13 pb0 = 2.9354831097821e-19   b1 = -1.91069189473616e-09 lb1 = 3.48786669964645e-15 wb1 = 1.45411716309218e-15 pb1 = -2.65441374640567e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.0975624497268945+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.35966435204754e-07 wvoff = -2.01948891952099e-07 pvoff = 3.83070697498373e-13   nfactor = {0.0885282131974474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.40403701136627e-06 wnfactor = 8.62108969723082e-07 pnfactor = 1.6583304412348e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.13819903971338 leta0 = -2.34666127187633e-06 weta0 = -9.30129612846585e-07 peta0 = 1.91852068438265e-12   etab = -0.464578826140316 letab = 9.57226610097737e-07 wetab = 3.58440198828912e-07 petab = -7.39332368270866e-13   dsub = -0.953068541985401 ldsub = 2.50212127130368e-06 wdsub = 6.80582643546282e-07 pdsub = -1.40379562271901e-12   voffl = 0.0   minv = 0.0   pclm = 1.54499878099653 lpclm = -2.16145824665687e-06 wpclm = -9.23141229315415e-07 ppclm = 1.67680303462735e-12   pdiblc1 = 0.422896399515241 lpdiblc1 = -6.78533637033179e-08 wpdiblc1 = -1.87593984980048e-08 ppdiblc1 = 3.86938481991278e-14   pdiblc2 = 0.000428309910268827 lpdiblc2 = -8.67569834851117e-10 wpdiblc2 = -1.62337843392791e-10 ppdiblc2 = 6.6025725576873e-16   pdiblcb = -2.1909393226472 lpdiblcb = 2.89779419126278e-06 wpdiblcb = 1.33442031490922e-06 ppdiblcb = -1.87172749695869e-12   drout = 0.118533961160854 ldrout = 9.10584627419096e-07 wdrout = 5.19118041139026e-08 pdrout = -1.07075259813891e-13   pscbe1 = 796411832.204736 lpscbe1 = 7.40109124488845 wpscbe1 = 2.730747112877 ppscbe1 = -5.63254276341038e-6   pscbe2 = 1.12733505466262e-08 lpscbe2 = -4.82454565772884e-15 wpscbe2 = -6.68702564140786e-16 ppscbe2 = 2.06653034379591e-21   pvag = 0.0   delta = 0.01   alpha0 = -1.03828228227482e-10 lalpha0 = 2.16595620787195e-16 walpha0 = 2.93258835065146e-18 palpha0 = -3.11627981975961e-24   alpha1 = -1.06283808041525e-10 lalpha1 = 2.1920501320963e-16 walpha1 = 1.06372205834572e-20 palpha1 = -1.13035148063168e-26   beta0 = -6.18145195509054 lbeta0 = 1.8938011697744e-05 wbeta0 = 2.21523956266197e-06 pbeta0 = -4.56923730104996e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.38662286987765e-09 lagidl = -2.94707064398043e-15 wagidl = -7.46250256056581e-16 pagidl = 1.99533118681403e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.32528579988031 lkt1 = -1.86074455760653e-07 wkt1 = -7.61968826001941e-08 pkt1 = 7.00886610579279e-14   kt2 = 0.0556219761979061 lkt2 = -1.39369313775648e-07 wkt2 = -6.21431929048911e-08 pkt2 = 7.54626340262706e-14   at = -48292.4883455517 lat = -0.0729020660645745 wat = 0.0299022077003358 pat = 8.13210568640139e-8   ute = 2.84911485768174 lute = -7.31566395717419e-06 wute = -2.60816265301252e-06 pute = 5.06980452701955e-12   ua1 = 2.81085929732118e-09 lua1 = -6.94974376808334e-15 wua1 = -2.18537667574537e-15 pua1 = 5.14367098739923e-21   ub1 = -5.17425309499604e-19 lub1 = 3.94084578701754e-24 wub1 = 1.17778547074228e-24 pub1 = -3.44414424228746e-30   uc1 = 1.90842565816185e-11 luc1 = 1.79272180564689e-16 wuc1 = 4.42279656865398e-17 puc1 = -1.60503140511121e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.86 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.967830807191816+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.47334923183026e-08 wvth0 = -6.35828054725181e-08 pvth0 = 7.15423764888282e-14   k1 = 0.291225418416654 lk1 = 7.90919236432371e-08 wk1 = 7.60494164114627e-08 pk1 = -9.68240386034326e-15   k2 = 0.018772444886922 lk2 = -6.75201650349346e-08 wk2 = 3.89790017954053e-09 pk2 = 3.82126178501322e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -384661.468380326 lvsat = 0.268063404316035 wvsat = 0.274671214217358 pvsat = -1.61503626775256e-7   ua = 1.64497750146726e-09 lua = 1.99785980230735e-16 wua = -1.46518127851975e-15 pua = -5.16773224677256e-22   ub = -8.83349319266785e-19 lub = -1.78062390990339e-25 wub = 8.34197091184632e-25 pub = 4.44734096686338e-31   uc = -1.9234617078362e-10 luc = 8.22115732466661e-17 wuc = 8.63142809253058e-17 puc = -3.81024969846161e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0163487176677751 lu0 = 5.75736020028689e-10 wu0 = -5.84315582990454e-09 pu0 = -1.46801696921702e-15   a0 = -2.95847764465984 la0 = 2.35240056577194e-06 wa0 = 2.41907931170503e-06 pa0 = -1.39842223439016e-12   keta = -0.195764595333149 lketa = 5.32454635509341e-08 wketa = 1.16346682411042e-07 pketa = -3.64414734340808e-14   a1 = 0.0   a2 = 3.1847390452944 la2 = -1.34174480696635e-06 wa2 = -1.81488704945675e-06 pa2 = 1.02112441973225e-12   ags = 3.09786275441824 lags = -2.48156158334121e-07 wags = -1.72559785505077e-06 pags = 3.95338070837548e-13   b0 = -3.72970048629149e-07 lb0 = 2.09926038135938e-13 wb0 = 2.83845946342834e-13 pb0 = -1.59762573900258e-19   b1 = -2.29018824329963e-08 lb1 = 2.57939034308422e-14 wb1 = 1.74292989909489e-14 pb1 = -1.96302490135957e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.379570414074611+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.89469230804493e-08 wvoff = 1.28337881488884e-07 pvoff = 3.20954211425932e-14   nfactor = {-4.69534016823042+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.67948331773748e-06 wnfactor = 5.10048220228905e-06 pnfactor = -2.84552601387263e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -2.82572068142676 leta0 = 1.86555045275659e-06 weta0 = 1.86025922569317e-06 peta0 = -1.04665253022555e-12   etab = 0.927102023866288 letab = -5.21626344991581e-07 wetab = -7.16880384535416e-07 petab = 4.03344145794238e-13   dsub = 2.55911637314918 ldsub = -1.2300598825451e-06 wdsub = -1.31366934863228e-06 pdsub = 7.15372325745632e-13   voffl = 0.0   minv = 0.0   pclm = -1.72989374687815 lpclm = 1.31856699937881e-06 wpclm = 1.38090583547184e-06 ppclm = -7.7156493020405e-13   pdiblc1 = 0.717966350127612 lpdiblc1 = -3.81405905882146e-07 wpdiblc1 = -6.10285097368622e-08 ppdiblc1 = 8.36106120277647e-14   pdiblc2 = -0.000147563254369685 lpdiblc2 = -2.55625126925976e-10 wpdiblc2 = 4.28803752552347e-12 ppdiblc2 = 4.83194262921454e-16   pdiblcb = 0.5360422 wpdiblcb = -4.2697679018084e-7   drout = 0.428186110040857 ldrout = 5.81536487237548e-07 wdrout = 2.91632585459347e-07 pdrout = -3.61811671461253e-13   pscbe1 = 807176335.590528 lpscbe1 = -4.03767910398346 wpscbe1 = -5.46149422575354 ppscbe1 = 3.07284418819007e-6   pscbe2 = -2.24286997322146e-08 lpscbe2 = 3.0988533646478e-14 wpscbe2 = 2.26924550854288e-14 ppscbe2 = -2.27579234986274e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 14.6608437318365 lbeta0 = -3.20980370642073e-06 wbeta0 = -4.49552879581423e-06 pbeta0 = 2.56188016586447e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -3.53051799583713e-09 lagidl = 2.278070091281e-15 wagidl = 2.52459043895567e-15 pagidl = -1.48038842765239e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.494280418604177 lkt1 = -6.49435210916234e-09 wkt1 = -1.9503890096781e-08 pkt1 = 9.84453289008638e-15   kt2 = -0.162858111126688 lkt2 = 9.27959292587844e-08 wkt2 = 6.7890266536327e-08 pkt2 = -6.27158612474267e-14   at = -318740.965638317 lat = 0.214486762948855 wat = 0.224030457795103 pat = -1.24966998560189e-7   ute = -7.83628955510095 lute = 4.03905281721639e-06 wute = 4.23953275638971e-06 pute = -2.20681682743682e-12   ua1 = -9.32105036972779e-09 lua1 = 5.94208445669024e-15 wua1 = 6.22845427761703e-15 pua1 = -3.79718550921989e-21   ub1 = 5.92615488841851e-18 lub1 = -2.90634738733777e-24 wub1 = -4.20612336182853e-24 pub1 = 2.27700187173791e-30   uc1 = 3.71736961300134e-10 luc1 = -1.95469984271985e-16 wuc1 = -2.27009647019816e-16 puc1 = 1.27724253779935e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.87 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.19782668703525+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.46709295250464e-08 wvth0 = 1.43073095933524e-07 pvth0 = -4.47300865664651e-14   k1 = 0.246158259331544 lk1 = 1.04448419896564e-07 wk1 = 1.32423550762278e-07 pk1 = -4.14006340632171e-14   k2 = -0.19651930879277 lk2 = 5.36111566719e-08 wk2 = 1.61622898445394e-07 pk2 = -5.0529459724171e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 26414.978949778 lvsat = 0.0367761741431193 wvsat = -0.0278526566017205 pvsat = 8.70779885464872e-9   ua = 6.47104661694388e-09 lua = -2.5155438947628e-15 wua = -5.3645595554442e-15 pua = 1.67716517029496e-21   ub = -4.41927116558865e-18 lub = 1.8113816047805e-24 wub = 3.65634031870511e-24 pub = -1.14311092455933e-30   uc = -1.0410808735264e-10 luc = 3.25654744612263e-17 wuc = 4.18447896265445e-17 puc = -1.30822713392636e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0336620594983614 lu0 = -9.1654080008487e-09 wu0 = -1.90223939161714e-08 pu0 = 5.94712318916398e-15   a0 = 1.73580869822328 la0 = -2.88783313615129e-07 wa0 = -1.49425154444283e-07 pa0 = 4.67159814351517e-14   keta = -0.215128987108101 lketa = 6.41406062104096e-08 wketa = 1.16078365057212e-07 pketa = -3.62905078947567e-14   a1 = 0.0   a2 = 1.14549842976048 la2 = -1.94390545523577e-7   ags = 5.45178929877987 lags = -1.57256468140066e-06 wags = -2.30219542053003e-06 pags = 7.19753771883668e-13   b0 = 3.156636613236e-10 lb0 = -9.86884557488876e-17 wb0 = -2.40233367273767e-16 pb0 = 7.5106079477736e-23   b1 = 5.16337364100239e-08 lb1 = -1.6142668083757e-14 wb1 = -3.92954523517047e-14 pb1 = 1.22852516323322e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.750383681072721+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.79686711836833e-07 wvoff = 4.17212760430944e-07 pvoff = -1.30436562995609e-13   nfactor = {1.85373211573062+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -5.27361396579085e-09 wnfactor = 9.67963658354963e-08 pnfactor = -3.02622222220783e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.409355e-05 letab = -3.95779542849e-11 wetab = 1.29246970711411e-26 petab = 4.62223186652937e-33   dsub = 0.0538379229831509 ldsub = 1.79504974099413e-07 wdsub = -9.49918769205568e-08 pdsub = 2.96980704166889e-14   voffl = 0.0   minv = 0.0   pclm = 0.584258857080582 lpclm = 1.65368065926809e-08 wpclm = 2.15406690166228e-08 ppclm = -6.73443168001885e-15   pdiblc1 = -0.487495902387309 lpdiblc1 = 2.96832964948343e-07 wpdiblc1 = 1.97094613465743e-07 ppdiblc1 = -6.16192657647031e-14   pdiblc2 = -0.0151950010085201 lpdiblc2 = 8.21063515619371e-09 wpdiblc2 = 1.94242750311496e-09 ppdiblc2 = -6.07276649718854e-16   pdiblcb = 1.4877650452944 lpdiblcb = -5.3547543823075e-07 wpdiblcb = -9.60933469095069e-07 ppdiblcb = 3.00424317910944e-13   drout = 2.74996328064118 ldrout = -7.24783576474678e-07 wdrout = -7.90912387374304e-07 pdrout = 2.47269266963928e-13   pscbe1 = 800088964.269279 lpscbe1 = -0.0500546785392544   pscbe2 = 6.1960005932288e-08 lpscbe2 = -1.64917589311864e-14 wpscbe2 = -3.99611438170876e-14 ppscbe2 = 1.24933720806866e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.53419290576835 lbeta0 = 2.37282861056593e-07 wbeta0 = 1.30099340980578e-07 pbeta0 = -4.0673997765485e-14   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.04161082855673e-09 lagidl = -2.9438332621832e-16 wagidl = -2.39831649037012e-16 pagidl = 7.49804870916333e-23   bgidl = 653150899.046399 lbgidl = 195.150484462332   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.498011030447117 lkt1 = -4.39536812307436e-09 wkt1 = -4.51638730474632e-09 pkt1 = 1.41199429418138e-15   kt2 = 0.0266627801067464 lkt2 = -1.3835725943013e-08 wkt2 = -9.80728698558428e-08 pkt2 = 3.0661305885991e-14   at = 57372.1951841752 lat = 0.00287120637000982 wat = 0.00432420061092781 pat = -1.35190943059926e-9   ute = -1.248076092906 lute = 3.32273571273947e-07 wute = 7.14021614211091e-07 pute = -2.23230289423727e-13   ua1 = 2.28743207298934e-09 lua1 = -5.89288887915242e-16 wua1 = -1.17128180547998e-15 pua1 = 3.6618720110165e-22   ub1 = 1.16273785908896e-18 lub1 = -2.26267956789854e-25 wub1 = -3.58091857258278e-25 pub1 = 1.11953122069514e-31   uc1 = 5.401768370832e-11 luc1 = -1.67090453662817e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.88 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.978057264371246+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.03734323778155e-09 wvth0 = -8.65022233032302e-08 pvth0 = 2.70438820890748e-14   k1 = -2.74321143825988 lk1 = 1.03903898341215e-06 wk1 = 1.08261172551904e-06 pk1 = -3.3846556464282e-13   k2 = 1.21176312579496 lk2 = -3.86671447112739e-07 wk2 = -4.18910404225226e-07 pk2 = 1.30967310956166e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -599704.170855863 lvsat = 0.232524812900055 wvsat = 0.466758579127344 pvsat = -1.45926468661214e-7   ua = 3.15983035151189e-09 lua = -1.48033186397067e-15 wua = -1.10067852005609e-15 pua = 3.44113931153295e-22   ub = -4.40049800406215e-18 lub = 1.80551240110718e-24 wub = 2.34588236833938e-24 pub = -7.33411971872887e-31   uc = -2.0420082383202e-12 luc = 6.55739619083645e-19 wuc = 1.13800680389117e-18 puc = -3.55784171154929e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00975803774095953 lu0 = -1.6921024466581e-09 wu0 = 1.59656224251644e-09 pu0 = -4.99146026375855e-16   a0 = 1.93720018971809 la0 = -3.51745946733087e-07 wa0 = -1.58139212619125e-06 pa0 = 4.94403271548182e-13   keta = 0.184791693752576 lketa = -6.08897956125108e-08 wketa = -2.46070349879336e-07 pketa = 7.69309420455758e-14   a1 = 0.0   a2 = -0.218272849934465 la2 = 2.31976179817691e-07 wa2 = 1.34534511617137e-07 pa2 = -4.20606006429587e-14   ags = -2.44893826583886 lags = 8.97502982946609e-07 pags = 2.01948391736579e-28   b0 = -4.7464696425673e-07 lb0 = 1.48392677611296e-13 wb0 = 3.61226369901263e-13 pb0 = -1.12933089833191e-19   b1 = -6.23096900818116e-08 lb1 = 1.94803768877974e-14 wb1 = 4.74203036211801e-14 pb1 = -1.48253888835185e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {1.26774812088445+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.51257978463453e-07 wvoff = -1.00024776194818e-06 pvoff = 3.12715459799956e-13   nfactor = {10.3591420101473+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -2.66438795253643e-06 wnfactor = -3.4868023969693e-06 pnfactor = 1.09010692778369e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.60302605655797 leta0 = -3.5336240270171e-08 weta0 = 6.49000812569598e-07 peta0 = -2.02902316040134e-13   etab = -0.545625515689248 letab = 1.70563730099055e-07 wetab = 4.98272061174247e-07 petab = -1.55778780661394e-13   dsub = 1.78915485048611 ldsub = -3.63021039481257e-07 wdsub = 6.20581338647701e-08 pdsub = -1.94017308552138e-14   voffl = 0.0   minv = 0.0   pclm = 0.727655757054981 lpclm = -2.82945134215151e-08 wpclm = -2.90579508177718e-08 ppclm = 9.0846196277665e-15   pdiblc1 = 1.69991270391659 lpdiblc1 = -3.87034086909295e-07 wpdiblc1 = -1.25142211596527e-07 ppdiblc1 = 3.91242107491151e-14   pdiblc2 = 0.0517796284238272 lpdiblc2 = -1.27281790402765e-08 wpdiblc2 = -7.89474387727761e-09 ppdiblc2 = 2.46819693630432e-15   pdiblcb = -0.0157261184236561 lpdiblcb = -6.54269677882649e-08 wpdiblcb = -5.54961449502257e-07 ppdiblcb = 1.73502037649487e-13   drout = -1.538265090594 ldrout = 6.15879565051547e-7   pscbe1 = 799682270.466854 lpscbe1 = 0.0770932584628099   pscbe2 = -7.2974330037405e-08 lpscbe2 = 2.56938419977064e-14 wpscbe2 = 6.20741779277965e-14 ppscbe2 = -1.94067468389904e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.98250225849324 lbeta0 = 7.22400321639388e-07 wbeta0 = 3.07958245438709e-06 pbeta0 = -9.62794499374674e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.40070446405048e-08 lagidl = -1.37270106223181e-14 wagidl = -3.3415113848708e-14 pagidl = 1.04468343634324e-20   bgidl = 2199791916.2286 lbgidl = -288.388269867479 wbgidl = 21.8553275877075 pbgidl = -6.83280590636553e-6   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 0.0752341222406692 lkt1 = -1.83613586169077e-07 wkt1 = -1.14552878397007e-07 pkt1 = 3.58135827962836e-14   kt2 = 0.337380461485714 lkt2 = -1.10977880413971e-07 wkt2 = 5.29395592033938e-23 pkt2 = 2.52435489670724e-29   at = 442705.2643898 lat = -0.117598553720298 wat = -0.266712845166987 pat = 8.33845704873166e-8   ute = 0.739069806217757 lute = -2.88983748336307e-07 wute = -6.21974769332592e-07 pute = 1.94452947934603e-13   ua1 = 1.42232089775527e-09 lua1 = -3.18822260312411e-16 wua1 = -1.11222852862211e-16 pua1 = 3.4772490273136e-23   ub1 = -2.06256945713866e-19 lub1 = 2.01731840994092e-25 wub1 = 4.9106776553136e-25 pub1 = -1.53526444080194e-31   uc1 = 2.26617492345528e-10 luc1 = -7.0670304339001e-17 wuc1 = -1.73003336597947e-16 puc1 = 5.40874171473088e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.89 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.707595428096791+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.96616622677425e-08 wvth0 = 1.13377345258634e-07 pvth0 = -2.14544966676385e-14   k1 = 2.76102110628785 lk1 = -2.96496992731817e-07 wk1 = -2.38652480711641e-06 pk1 = 5.03278785362778e-13   k2 = -0.862060721021584 lk2 = 1.16517023431134e-07 wk2 = 9.94839943393683e-07 pk2 = -2.12062245889391e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2383811.70962028 lvsat = -0.491389513306915 wvsat = -1.1239218879846 pvsat = 2.40033058517894e-7   ua = -4.02742940620106e-09 lua = 2.63570469121281e-16 wua = -1.21472889947219e-15 pua = 3.71786887114059e-22   ub = 2.58078524006969e-18 lub = 1.11587797317518e-25 wub = 1.72892988300295e-24 pub = -5.83715854735825e-31   uc = 4.0322971490355e-12 luc = -8.18117691493566e-19 wuc = -2.49127536664197e-18 puc = 5.24817596138893e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00252938593216812 lu0 = 1.28929345854224e-09 wu0 = -2.69210473491985e-09 pu0 = 5.41447551695331e-16   a0 = -3.26579179983514 la0 = 9.10697623628133e-07 wa0 = 3.52700930252263e-06 pa0 = -7.45089034312099e-13   keta = -3.14447583421041 lketa = 7.46917018837373e-07 wketa = 2.03876156925514e-06 pketa = -4.77456105149375e-13   a1 = 0.0   a2 = -1.11722629815691 la2 = 4.5009644658749e-07 wa2 = -3.13913860439986e-07 pa2 = 6.6750015456238e-14   ags = 19.3498474922719 lags = -4.39171079582987e-06 wags = -1.01547782567287e-05 pags = 2.46393508665614e-12   b0 = -9.69285283192636e-07 lb0 = 2.68410730041266e-13 wb0 = 7.37667004348547e-13 pb0 = -2.04271892494211e-19   b1 = 6.68773396242748e-07 lb1 = -1.57908161011821e-13 wb1 = -5.08964776778053e-13 pb1 = 1.20174774254391e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-6.80565782361187+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.50765709309725e-06 wvoff = 5.05965327601729e-06 pvoff = -1.15764680824991e-12   nfactor = {-21.9203242483037+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.1678371814816e-06 wnfactor = 1.72150213306424e-05 pnfactor = -3.93294217783656e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.208617739578622 leta0 = 1.6159938713682e-07 weta0 = -7.06421550433318e-07 peta0 = 1.25974655274168e-13   etab = 2.39212151265688 letab = -5.42245333364792e-07 wetab = -1.79080382272017e-06 petab = 3.9963801365498e-13   dsub = 0.622365523453393 ldsub = -7.99136107486921e-08 wdsub = -2.17378608918663e-07 pdsub = 4.84002415402726e-14   voffl = 0.0   minv = 0.0   pclm = 1.67424949550111 lpclm = -2.57974124930606e-07 wpclm = 1.01560694170476e-06 ppclm = -2.44390780564115e-13   pdiblc1 = 0.515568993053107 lpdiblc1 = -9.96672975928012e-08 wpdiblc1 = 4.39534666129748e-07 ppdiblc1 = -9.7887857508633e-14   pdiblc2 = -0.0128051402316259 lpdiblc2 = 2.94254005674533e-09 wpdiblc2 = 2.16744307974397e-08 ppdiblc2 = -4.70640846841975e-15   pdiblcb = -2.42980992756405 lpdiblcb = 5.20321499493941e-07 wpdiblcb = 1.38767519428466e-06 ppdiblcb = -2.97855432325683e-13   drout = 1.0   pscbe1 = 1634204399.62469 lpscbe1 = -202.409687116136 wpscbe1 = -467.893796057275 ppscbe1 = 0.000113528814887745   pscbe2 = 2.085092045711e-07 lpscbe2 = -4.26047598726319e-14 wpscbe2 = -1.48373665034095e-13 ppscbe2 = 3.1655896881597e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 38.0182900152037 lbeta0 = -6.80806114807334e-06 wbeta0 = -1.39804776230218e-05 pbeta0 = 3.17662435768768e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -7.33418209152674e-08 lagidl = 1.47462834184033e-14 wagidl = 5.52376032971018e-14 pagidl = -1.10636836193926e-20   bgidl = 1090894703.41325 lbgidl = -19.3276679443879 wbgidl = -50.9957643713169 pbgidl = 1.08436373443886e-5   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.481232744561552 lkt1 = -4.85935785419207e-08 wkt1 = 2.67290049593018e-07 pkt1 = -5.683602156536e-14   kt2 = -0.12   at = -77498.6682373276 lat = 0.0086226880844828 wat = 0.309159856765644 pat = -5.63440301642132e-8   ute = -1.53576181598151 lute = 2.62976846810878e-07 wute = 9.84152242070662e-07 pute = -1.9525449785826e-13   ua1 = 1.44639081629341e-09 lua1 = -3.24662537206668e-16 wua1 = -7.54923599526532e-16 pua1 = 1.90958752042273e-22   ub1 = 2.44139278733235e-18 lub1 = -4.40688594932776e-25 wub1 = -1.14582478623984e-24 pub1 = 2.43645890896467e-31   uc1 = -5.79236678308897e-10 luc1 = 1.24860539920247e-16 wuc1 = 4.03674452061875e-16 puc1 = -8.5836528137533e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.90 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0379169+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47866595   k2 = 0.0148198355   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24491.02   ua = -9.0151189e-10   ub = 7.0651505e-19   uc = -6.8009552e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0066877133   a0 = 1.2509318   keta = 0.0074076058   a1 = 0.0   a2 = 0.8   ags = 0.23496304   b0 = -3.2678e-8   b1 = 1.9071e-9   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.19048746+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.3892827+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00083787503   pdiblcb = -0.225   drout = 0.56   pscbe1 = 790097310.0   pscbe2 = 9.5178184e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1731672e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.52561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.91 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0379169+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47866595   k2 = 0.0148198355   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 24491.02   ua = -9.0151189e-10   ub = 7.0651505e-19   uc = -6.8009552e-11   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0066877133   a0 = 1.2509318   keta = 0.0074076058   a1 = 0.0   a2 = 0.8   ags = 0.23496304   b0 = -3.2678e-8   b1 = 1.9071e-9   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.19048746+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}   nfactor = {1.3892827+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.0017402344   pdiblc1 = 0.39   pdiblc2 = 0.00083787503   pdiblcb = -0.225   drout = 0.56   pscbe1 = 790097310.0   pscbe2 = 9.5178184e-9   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.1731672e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.52561   kt2 = -0.052484   at = 10000.0   ute = -1.2595   ua1 = -2.5605e-10   ub1 = 4.9434e-19   uc1 = 8.1951e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.92 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.0545024165031+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.33723015607515e-7   k1 = 0.495199413953725 lk1 = -1.33303334744933e-7   k2 = 0.0077526009474457 lk2 = 5.6980553858337e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -7466.68585431 lvsat = 0.257663413613782   ua = -9.5079223739613e-10 lua = 3.97329601569238e-16   ub = 8.01070674372721e-19 lub = -7.62367770181221e-25   uc = -6.32636666507766e-11 luc = -3.82643555602928e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00629912532697635 lu0 = 3.13304415764345e-9   a0 = 1.2539489181107 la0 = -2.43259311298079e-8   keta = 0.0041253241822056 lketa = 2.64638484983306e-8   a1 = 0.0   a2 = 0.8   ags = 0.235899528841975 lags = -7.55057052388457e-9   b0 = -3.5828575769e-08 lb0 = 2.54019519170187e-14   b1 = 3.67664292047e-09 lb1 = -1.42671839932124e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.200872629170475+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 8.37318595902992e-8   nfactor = {0.884435637253649+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.0703991122871e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -0.402583092873373 lpclm = 3.25991262276074e-06 wpclm = 9.26442286059391e-23 ppclm = -1.38839519318898e-28   pdiblc1 = 0.39   pdiblc2 = 0.00125213717903229 lpdiblc2 = -3.34004574474937e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 780039548.825947 lpscbe1 = 81.0920874368603   pscbe2 = 9.45533705887899e-09 lpscbe2 = 5.03764435213175e-16   pvag = 0.0   delta = 0.01   alpha0 = 1.79950418418211e-10 lalpha0 = -6.44611281654569e-16   alpha1 = 2.0156591584996e-10 lalpha1 = -8.18889212636695e-16   beta0 = -17.9894678937345 lbeta0 = 0.000169230481439804   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.2631396617684e-09 lagidl = -8.78805338920745e-15   bgidl = 673331505.26195 lbgidl = 2633.8098190778   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.660347389269999 lkt1 = 1.08633879474909e-06 wkt1 = 4.2351647362715e-22   kt2 = -0.046345693212273 lkt2 = -4.94909455623856e-8   at = -43627.8504630735 lat = 0.432381945001894   ute = -2.169175431175 lute = 7.33438369905793e-6   ua1 = -8.9668738622e-10 lua1 = 5.16522733435805e-15 pua1 = 1.50463276905253e-36   ub1 = 5.6646681563422e-19 lub1 = -5.81532404551458e-25   uc1 = 6.16128714520936e-11 luc1 = -4.30688153984964e-16 wuc1 = 6.16297582203915e-33 puc1 = 7.05296610493373e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.93 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.9884442200884+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.34647523358303e-7   k1 = 0.47574838516156 lk1 = -5.42808460347892e-8   k2 = 0.028963061019078 lk2 = -2.91898672261589e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 80360.830639533 lvsat = -0.0991479923397309   ua = -1.18417577807895e-09 lua = 1.34548244252181e-15   ub = 8.20404075558569e-19 lub = -8.40912380508097e-25   uc = -7.91412024139669e-11 luc = 2.62403245776042e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00565267952897999 lu0 = 5.75931942152376e-9   a0 = 1.3368208826228 la0 = -3.61004723291323e-7   keta = 0.0270829359938964 lketa = -6.68046176370933e-8   a1 = 0.0   a2 = 0.8   ags = -0.11320416886595 lags = 1.41073137772485e-06 pags = 4.03896783473158e-28   b0 = -5.987189287253e-08 lb0 = 1.2308124562787e-13   b1 = 2.54064563285e-10 lb1 = -3.62487101335046e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1689708076647+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.58736927282786e-8   nfactor = {1.379840487444+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.05774854251948e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.1619898605 leta0 = -3.33095122881999e-7   etab = -0.1416766705 letab = 2.91196365286779e-7   dsub = 0.8693957 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = 0.50209638586452 lpclm = -4.15472605380022e-7   pdiblc1 = 0.39   pdiblc2 = 0.000575520296916849 lpdiblc2 = -5.91196288025677e-10   pdiblcb = -0.4312638 lpdiblcb = 8.379751519044e-7   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.63207382525211e-09 lpscbe2 = -2.14253067851319e-16   pvag = 0.0   delta = 0.01   alpha0 = 3.93997587660097e-11 lalpha0 = -7.36048308264681e-17   alpha1 = 5.92445188998808e-16 lalpha1 = -2.27029018019908e-21 walpha1 = 9.4039548065783e-38 palpha1 = -4.48415508583941e-43   beta0 = 44.978935787469 lbeta0 = -8.65873481547934e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.5984741217841e-10 lagidl = 1.05566597091767e-15 pagidl = -1.88079096131566e-37   bgidl = 1653336989.4761 lbgidl = -1347.597701299 wbgidl = -9.09494701772928e-13   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.292092426537939 lkt1 = -4.09747810534757e-7   kt2 = -0.059587033782843 lkt2 = 4.30382781055369e-9   at = 86384.839460565 lat = -0.0958125495640969   ute = 0.256564572347719 lute = -2.5205198173736e-06 pute = 8.07793566946316e-28   ua1 = 7.70305797178011e-10 lua1 = -1.60716251825568e-15   ub1 = 3.2750382410512e-19 lub1 = 3.89287725428343e-25   uc1 = -1.37767291420899e-10 luc1 = 3.79321272149044e-16 puc1 = -9.4039548065783e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.94 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.087351210829+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.93617942089061e-8   k1 = 0.4116737627374 lk1 = 7.78819050129338e-8   k2 = 0.00262944467909798 lk2 = 2.51268505141047e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -25075.666742956 lvsat = 0.118329333748291   ua = 6.51366217055801e-10 lua = -2.44057622723894e-15 pua = -7.52316384526264e-37   ub = -4.0467067035072e-19 lub = 1.68597334324475e-24   uc = -1.1038572076075e-10 luc = 9.06864554113759e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0131540234289 lu0 = -9.71323755751944e-9   a0 = 1.0984667752 la0 = 1.30633516135022e-7   keta = -0.0115733216886196 lketa = 1.29292483966562e-8   a1 = 0.0   a2 = 1.2250552 la2 = -8.767350076176e-7   ags = 0.697188575545621 lags = -2.60815491822746e-07 wags = -4.2351647362715e-22   b0 = -6.686273779694e-08 lb0 = 1.37500828021065e-13 wb0 = -4.53595020502082e-30 pb0 = -4.13774011489445e-36   b1 = 6.8112234507e-10 lb1 = -1.24335271024049e-15 wb1 = 9.86076131526265e-32   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.262390673143539+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.46817671763265e-7   nfactor = {1.6251487556862+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.55176638672893e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.519661301 leta0 = 1.07290446557204e-06 weta0 = 8.31316515615793e-23 peta0 = -3.94430452610506e-31   etab = 0.174303951 letab = -3.60557271882738e-07 wetab = 2.27474668452083e-23 petab = 3.94430452610506e-31   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = -0.10040548505586 lpclm = 8.27270648651448e-7   pdiblc1 = 0.389459701708899 lpdiblc1 = 1.11443978655844e-9   pdiblc2 = 0.0001389594061663 lpdiblc2 = 3.09270794550254e-10   pdiblcb = 0.1875276 lpdiblcb = -4.383675038088e-7   drout = 0.21106141117068 ldrout = 7.19733992985731e-7   pscbe1 = 801279107.986979 lpscbe1 = -2.63833674004854   pscbe2 = 1.00814570239272e-08 lpscbe2 = -1.14116793000014e-15   pvag = 0.0   delta = 0.01   alpha0 = -9.86011912048635e-11 lalpha0 = 2.11041172619554e-16 walpha0 = 9.24446373305873e-33 palpha0 = -1.46936793852786e-38   alpha1 = -1.06264848290221e-10 lalpha1 = 2.19184865857423e-16 walpha1 = 1.83700614773623e-32 palpha1 = 2.23303748626666e-38   beta0 = -2.2330153443294 lbeta0 = 1.07938163037969e-05 pbeta0 = 3.23117426778526e-27   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.65085646496596e-11 lagidl = 6.09401911584975e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.461098903779081 lkt1 = -6.11486283310467e-8   kt2 = -0.0551418716996158 lkt2 = -4.86493241846932e-9   at = 5005.12046236999 lat = 0.072044351270902   ute = -1.79966673666628 lute = 1.72074101738842e-6   ua1 = -1.08434978988362e-09 lua1 = 2.21832057252995e-15 wua1 = -5.54667823983524e-32 pua1 = 2.35098870164458e-38   ub1 = 1.58185611842556e-18 lub1 = -2.19798698222418e-24   uc1 = 9.79160551282162e-11 luc1 = -1.0680815441033e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.95 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.08116061638+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.27834333048099e-8   k1 = 0.426775679005719 lk1 = 6.18340349134001e-8   k2 = 0.0257200509307108 lk2 = 5.89894868103335e-10   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 104911.71206378 lvsat = -0.019800194492141   ua = -9.66557385783196e-10 lua = -7.21309125765311e-16   ub = 6.03521171374798e-19 lub = 6.14630380937224e-25   uc = -3.849984527494e-11 luc = 1.42977924568857e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00593389356023999 lu0 = -2.04085319414632e-9   a0 = 1.3532823472 la0 = -1.40143193663914e-07 wa0 = -8.470329472543e-22   keta = 0.0116113960112492 lketa = -1.1707713650497e-08 wketa = 2.8951321439356e-24 pketa = -1.97215226305253e-30   a1 = 0.0   a2 = -0.0501104000000003 la2 = 4.783044152352e-7   ags = 0.0221621118448798 lags = 4.5649327951128e-7   b0 = 1.32956147908e-07 lb0 = -7.48343130466612e-14   b1 = 8.16404984616e-09 lb1 = -9.19499582414377e-15 wb1 = -7.88860905221012e-31 pb1 = -1.1284745767894e-36   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.15082134406012+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.82598630447178e-8   nfactor = {4.3957446063+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.39237404677562e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = -0.350663507025 letab = 1.97293097778032e-7   dsub = 0.21763591297652 ldsub = 4.50176887064566e-8   voffl = 0.0   minv = 0.0   pclm = 0.731428833619079 lpclm = -5.6668108076652e-8   pdiblc1 = 0.60918931029556 lpdiblc1 = -2.32378592022753e-7   pdiblc2 = -0.00013992026864504 lpdiblc2 = 6.05618934432429e-10 ppdiblc2 = -1.97215226305253e-31   pdiblcb = -0.225   drout = 0.947991189693241 ldrout = -6.33555930039246e-8   pscbe1 = 797441784.026039 lpscbe1 = 1.43934951915708   pscbe2 = 1.80182667979836e-08 lpscbe2 = -9.57512359468389e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.64802616514679 lbeta0 = 1.35648411625014e-6   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 9.69304725084159e-10 lagidl = -3.60569974746822e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.529044096090081 lkt1 = 1.105251493593e-8   kt2 = -0.0418506957552119 lkt2 = -1.8988641041679e-8   at = 80570.2765375879 lat = -0.00825405505055543   ute = -0.279758591138324 lute = 1.05628865440884e-7   ua1 = 1.7805285803352e-09 lua1 = -8.26008049042636e-16 wua1 = -7.88860905221012e-31   ub1 = -1.57082726698536e-18 lub1 = 1.15217418508211e-24 wub1 = -3.67341984631965e-40   uc1 = -3.28843791619844e-11 luc1 = 3.21853574829406e-17 wuc1 = -3.08148791101958e-33 puc1 = 2.93873587705572e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.96 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.94281361327088+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.50558478304985e-8   k1 = 0.482189614481439 lk1 = 3.06560490852116e-8   k2 = 0.0915568794964424 lk2 = -3.64524066824627e-08 pk2 = 6.31088724176809e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -23229.51588808 lvsat = 0.0522969297202376   ua = -3.0907288706116e-09 lua = 4.7383047011557e-16   ub = 2.097779278576e-18 lub = -2.26096011982243e-25   uc = -2.95240549455508e-11 luc = 9.2476717375388e-18   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.000243400583200007 lu0 = 1.43472722813048e-9   a0 = 1.46947373368 la0 = -2.05516882970247e-07 wa0 = -8.470329472543e-22   keta = -0.00823124384170799 lketa = -5.43490448908891e-10   a1 = 0.0   a2 = 1.14549842976048 la2 = -1.94390545523577e-7   ags = 1.34836281761672 lags = -2.89677633182776e-7   b0 = -1.125276e-10 lb0 = 3.51804038088e-17   b1 = -1.84063645872e-08 lb1 = 5.75452901181303e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.00674485955279969+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.28030420455117e-8   nfactor = {2.0262616791672+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -5.9212911619476e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 6.409355e-05 letab = -3.95779542849e-11 wetab = -6.46234853557053e-27 petab = 1.23259516440783e-32   dsub = -0.115475324613119 ldsub = 2.32438729201417e-7   voffl = 0.0   minv = 0.0   pclm = 0.622652883441919 lpclm = 4.53337497912547e-9   pdiblc1 = -0.13619503149784 lpdiblc1 = 1.87002963275202e-07 ppdiblc1 = 5.04870979341448e-29   pdiblc2 = -0.0117328238262779 lpdiblc2 = 7.12822700629187e-09 wpdiblc2 = -8.27180612553028e-25 ppdiblc2 = -1.18329135783152e-30   pdiblcb = -0.225   drout = 1.34024332129712 ldrout = -2.84051547825269e-7   pscbe1 = 800088964.269278 lpscbe1 = -0.0500546785397091   pscbe2 = -9.2666216138888e-09 lpscbe2 = 5.77639145159516e-15 wpscbe2 = -7.88860905221012e-31 ppscbe2 = 3.76158192263132e-37   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.76608159610321 lbeta0 = 1.64785644687687e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 6.1413558866032e-10 lagidl = -1.60738322167585e-16   bgidl = 653150899.046398 lbgidl = 195.150484462331   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.506061026159999 lkt1 = -1.87863356338981e-9   kt2 = -0.148142020416 lkt2 = 4.08148972828174e-8   at = 65079.637888 lat = 0.000461566897971444   ute = 0.0245939740000001 lute = -6.5611453103412e-8   ua1 = 1.9974275928e-10 lua1 = 6.34021237442192e-17   ub1 = 5.2447596496e-19 lub1 = -2.67230347331647e-26   uc1 = 5.401768370832e-11 luc1 = -1.67090453662817e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.97 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.13223857783257+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 4.41655942401396e-8   k1 = -0.813567419469425 lk1 = 4.35758936665543e-7   k2 = 0.4650984288698 lk2 = -1.53235689595451e-07 wk2 = 5.29395592033938e-23 pk2 = -2.52435489670724e-29   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 232244.975086 lvsat = -0.0275741041889168   ua = 1.19798413021857e-09 lua = -8.66984185037976e-16   ub = -2.19204033057143e-19 lub = 4.98281016600118e-25   uc = -1.36281915230571e-14 luc = 2.15909380130796e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0126037456797143 lu0 = -2.58177888521451e-9   a0 = -0.881468577428571 la0 = 5.29477019290113e-7   keta = -0.253803388541297 lketa = 7.62316937256813e-08 wketa = -2.64697796016969e-23 pketa = 6.31088724176809e-30   a1 = 0.0   a2 = 0.0215210757580024 la2 = 1.5700748647705e-7   ags = -2.44893826583885 lags = 8.97502982946609e-7   b0 = 1.69201876171429e-07 lb0 = -5.28989361624831e-14   b1 = 2.22121223971429e-08 lb1 = -6.94435352199795e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.515090606662572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.06125155639393e-7   nfactor = {4.14427546896858+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -7.21384506835397e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.75980323404943 leta0 = -3.96988743486745e-07 peta0 = -2.01948391736579e-28   etab = 0.342493169811142 letab = -1.07095919498416e-07 wetab = 5.4697318005069e-23 petab = 9.86076131526265e-30   dsub = 1.89976708939571 ldsub = -3.97602628629478e-7   voffl = 0.0   minv = 0.0   pclm = 0.675862949280855 lpclm = -1.21021135846287e-8   pdiblc1 = 1.47685958670629 lpdiblc1 = -3.172992064509e-7   pdiblc2 = 0.0377080596946343 lpdiblc2 = -8.32887193591908e-9   pdiblcb = -1.00488780626506 lpdiblcb = 2.43822563975097e-7   drout = -1.538265090594 ldrout = 6.15879565051547e-7   pscbe1 = 799682270.466858 lpscbe1 = 0.0770932584628099   pscbe2 = 3.76665057638886e-08 lpscbe2 = -8.89668762553839e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 12.47154114788 lbeta0 = -9.93681818660703e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.55519579598486e-08 lagidl = 4.89339683265114e-15 wagidl = -2.36658271566304e-30 pagidl = 1.1284745767894e-36   bgidl = 2238746789.12 lbgidl = -300.567043418498   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.128944597999999 lkt1 = -1.19779559430476e-7   kt2 = 0.337380461485714 lkt2 = -1.10977880413971e-07 wkt2 = 5.29395592033938e-23   at = -32682.9419999998 lat = 0.031025864348996   ute = -0.369536229714286 lute = 5.76086255254147e-8   ua1 = 1.22407760542857e-09 lua1 = -2.56843873885978e-16   ub1 = 6.69020824e-19 lub1 = -7.19132503737123e-26   uc1 = -8.17431561011428e-11 luc1 = 2.57349520700691e-17 wuc1 = 1.07852076885685e-32 puc1 = 1.10202595389589e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.98 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.16414265538985+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.13023755426483e-07 wvth0 = -9.36746706924495e-07 pvth0 = 2.27290347474746e-13   k1 = -5.48591798200817 lk1 = 1.56944873245882e-06 wk1 = 2.24035604224718e-06 pk1 = -5.43595509378773e-13   k2 = 2.84425737771021 lk2 = -7.30510058624189e-07 wk2 = -1.08456091661862e-06 pk2 = 2.63155691686508e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 798655.073847516 lvsat = -0.165006717732214 wvsat = -0.234582121706052 pvsat = 5.69185368465129e-8   ua = -2.95149347116528e-08 lua = 6.58513701691602e-15 wua = 1.30848371496101e-14 pua = -3.1748787163071e-21   ub = 3.1025012163808e-17 lub = -7.08275311297484e-24 wub = -1.42294817675904e-23 pub = 3.4526129971246e-30   uc = 1.25243887305262e-13 luc = -1.21047054496664e-20 wuc = -2.99253609163667e-19 puc = 7.2610297220254e-26   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.064726244214353 lu0 = 1.61814152027022e-08 wu0 = 3.22029574688054e-08 pu0 = -7.813661194316e-15   a0 = -12.2812038187683 la0 = 3.2954859787783e-06 wa0 = 8.58503589553132e-06 pa0 = -2.08305593961993e-12   keta = -0.432034455886139 lketa = 1.19477323444099e-07 wketa = 5.16967490989056e-07 pketa = -1.25435958078603e-13   a1 = 0.0   a2 = -9.0775652836831 la2 = 2.36479160255912e-06 wa2 = 4.15217223674539e-06 pa2 = -1.00747476717943e-12   ags = 24.4355257693518 lags = -5.62568960162398e-06 wags = -1.30080583857938e-05 pags = 3.15624927061224e-12   b0 = -1.48853757152547e-06 lb0 = 3.49331647947798e-13 wb0 = 1.02898945054984e-12 pb0 = -2.49671942302511e-19   b1 = -1.28073987058189e-06 lb1 = 3.09201312150449e-13 wb1 = 5.84794435370431e-13 pb1 = -1.41893352209411e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {12.3665216329514+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.01944347495605e-06 wvoff = -5.69674846508775e-06 pvoff = 1.38224765407196e-12   nfactor = {68.4183685934935+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.63167219143839e-05 wnfactor = -3.34687976464437e-05 pnfactor = 8.12080212333782e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -7.72042519324649 leta0 = 1.90327492165548e-06 weta0 = 3.5080194293489e-06 peta0 = -8.5117881829836e-13   etab = -1.62729796214823 letab = 3.70850261177942e-07 wetab = 4.64260122147331e-07 petab = -1.12647147517584e-13   dsub = 0.0569851637544083 ldsub = 4.95262922442782e-08 wdsub = 9.98236319236481e-08 pdsub = -2.42210064026902e-14   voffl = 0.0   minv = 0.0   pclm = 18.1309947193706 lpclm = -4.24738037601567e-06 wpclm = -8.21732160353449e-06 ppclm = 1.9938344792384e-12   pdiblc1 = 7.53649800604412 lpdiblc1 = -1.78759775324219e-06 wpdiblc1 = -3.49950279336256e-06 ppdiblc1 = 8.49112358775904e-13   pdiblc2 = 0.152679283588389 lpdiblc2 = -3.62252597590519e-08 wpdiblc2 = -7.11693144082737e-08 ppdiblc2 = 1.72683801093947e-14   pdiblcb = -2.51035948308532 lpdiblcb = 6.09107200695411e-07 wpdiblcb = 1.43286689412333e-06 ppdiblcb = -3.47667957456298e-13   drout = 1.0   pscbe1 = 801445283.976006 lpscbe1 = -0.350680813367944 wpscbe1 = -0.680789743677451 ppscbe1 = 1.65185461826339e-7   pscbe2 = -4.23438065912289e-08 lpscbe2 = 1.05168545436826e-14 wpscbe2 = -7.63453977495752e-15 ppscbe2 = 1.85242946191615e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 14.9689444110145 lbeta0 = -1.59964675162111e-06 wbeta0 = -1.04882205668715e-06 pbeta0 = 2.54484086190452e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 1.73223637632492e-08 lagidl = -3.08316284159784e-15 wagidl = 4.37116966386056e-15 pagidl = -1.06061186489981e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = 2.49514039988792 lkt1 = -7.56482295148005e-07 wkt1 = -1.40258088738983e-06 pkt1 = 3.40319421354494e-13   kt2 = -0.12   at = 1098628.74400839 lat = -0.243473340520708 wat = -0.350697254081001 pat = 8.50924803357061e-8   ute = 6.95369079722695 lute = -1.71928453383755e-06 wute = -3.77878892883956e-06 pute = 9.16877788115774e-13   ua1 = -7.69845695024031e-10 lua1 = 2.26957687889242e-16 wua1 = 4.8847860850333e-16 pua1 = -1.18523472610031e-22   ub1 = 5.37449209124823e-19 lub1 = -3.99889768836298e-26 wub1 = -7.76320924464173e-26 pub1 = 1.88364956470143e-32   uc1 = 7.58416166831534e-10 luc1 = -1.7811962572767e-16 wuc1 = -3.46805243011972e-16 puc1 = 8.41481305539389e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.99 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.02634743687523+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -5.44970536311051e-9   k1 = 0.5331222043272 wk1 = -2.56511938420438e-8   k2 = -0.0486465635545884 wk2 = 2.98953522367513e-8   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -174004.013986969 wvsat = 0.0934995374982968   ua = -1.29760299696875e-09 wua = 1.86575626426997e-16   ub = 1.13848463589725e-18 wub = -2.03475904074128e-25   uc = -2.21696422835493e-11 wuc = -2.15925319206383e-17   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00536780967883877 wu0 = 6.21730305499754e-10   a0 = 0.348643534644155 wa0 = 4.25015849547401e-7   keta = -0.0379454693240326 wketa = 2.13632122831896e-8   a1 = 0.0   a2 = 0.276631393076923 wa2 = 2.46528700015981e-7   ags = 0.494527949826646 wags = -1.22266026167545e-7   b0 = 7.05922015615385e-08 wb0 = -4.86446229379905e-14   b1 = -1.83885836621538e-08 wb1 = 9.560123482725e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.249015312216938+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 2.75690882695416e-8   nfactor = {2.34285899011308+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -4.49174673562702e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.00593665147881314 wpclm = -1.97668953292171e-9   pdiblc1 = 0.39   pdiblc2 = -0.00330061165006257 wpdiblc2 = 1.94940187044737e-9   pdiblcb = -0.225   drout = 0.56   pscbe1 = 1170341077.89128 wpscbe1 = -179.110860963796   pscbe2 = 8.51699517285954e-09 wpscbe2 = 4.71429974723342e-16   pvag = 0.0   delta = 0.01   alpha0 = 3.62340153846154e-10 walpha0 = -1.23573283216031e-16   alpha1 = 3.62340153846154e-10 walpha1 = -1.23573283216031e-16   beta0 = -67.8318415384615 wbeta0 = 3.33647864683283e-5   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 2.77148754691129e-09 wagidl = -7.52876332513858e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.01642219383077 wkt1 = 2.31193255568872e-7   kt2 = -0.0355196086772415 wkt2 = -7.99094421033305e-9   at = -186853.8208675 wat = 0.0927264568598331   ute = -3.77471245901538 wute = 1.18477121016202e-6   ua1 = -2.55288928195512e-09 wua1 = 1.08190822841856e-15   ub1 = 1.14831103222126e-18 wub1 = -3.08047953753774e-25   uc1 = -1.51790770957345e-10 wuc1 = 7.53600966246637e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.100 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.10528021361434+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.5835997260516e-06 wvth0 = 3.1730963444189e-08 pvth0 = -7.45942298878738e-13   k1 = 0.551249371125776 lk1 = -3.63678785445444e-07 wk1 = -3.41898543706117e-08 pk1 = 1.71308055189549e-13   k2 = -0.0979475546729789 lk2 = 9.89107937849482e-07 wk2 = 5.31181995553384e-08 pk2 = -4.65911579082083e-13   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -277584.024542017 lvsat = 2.0780882558021 wvsat = 0.14229009354617 pvsat = -9.78867263807186e-7   ua = -1.32556823713085e-09 lua = 5.6105648995519e-16 wua = 1.99748434676479e-16 pua = -2.64281283352773e-22   ub = 1.2485268992687e-18 lub = -2.20773809472223e-24 wub = -2.55310453905599e-25 pub = 1.03993780916177e-30   uc = -1.40762904591584e-11 luc = -1.62373987859393e-16 wuc = -2.54048421693734e-17 puc = 7.64850004640616e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00659242038892644 lu0 = -2.45689213674119e-08 wu0 = 4.48869824764932e-11 pu0 = 1.15729987725327e-14   a0 = -0.228691719993713 la0 = 1.15828682184374e-05 wa0 = 6.96965118029584e-07 pa0 = -5.45601972792282e-12   keta = -0.0637795176399231 lketa = 5.18299159436221e-07 wketa = 3.3532139236813e-08 pketa = -2.44140776318988e-13   a1 = 0.0   a2 = -0.0750129084384978 la2 = 7.05491232606676e-06 wa2 = 4.12168005419269e-07 pa2 = -3.3231614228776e-12   ags = 0.651746195769587 lags = -3.15421275534818e-06 wags = -1.96322454616649e-07 pags = 1.48576731554727e-12   b0 = 1.98458530207319e-07 lb0 = -2.56533586400933e-12 wb0 = -1.08875059689222e-13 pb0 = 1.20838144912185e-18   b1 = -3.47728814437098e-08 lb1 = 3.28712235275561e-13 wb1 = 1.72778191552043e-14 pb1 = -1.54837334471118e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.309514260124503+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.21376849125032e-06 wvoff = 5.6066645789606e-08 pvoff = -5.7173618040923e-13   nfactor = {3.78099376049076+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.88527772933006e-05 wnfactor = -1.1265968396979e-06 pnfactor = 1.35908756923464e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.18685961114232e-06 lcit = 1.76814845264831e-10 wcit = 4.15136103767638e-12 pcit = -8.32872537062056e-17   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 1.08607158538335 lpclm = -2.16703561700807e-05 wpclm = -5.1076582509617e-07 ppclm = 1.02076522451384e-11   pdiblc1 = 0.39   pdiblc2 = -0.00667915420608639 lpdiblc2 = 6.77824762691007e-08 wpdiblc2 = 3.54083798883046e-09 ppdiblc2 = -3.1928406743245e-14   pdiblcb = -0.225   drout = 0.56   pscbe1 = 1421313828.56394 lpscbe1 = -5035.17544460989 wpscbe1 = -297.329617580699 ppscbe1 = 0.00237178011881502   pscbe2 = 7.78835310382083e-09 lpscbe2 = 1.46184820626945e-14 wpscbe2 = 8.14651137935886e-16 ppscbe2 = -6.88592195147215e-21   pvag = 0.0   delta = 0.01   alpha0 = 5.38602961623308e-10 lalpha0 = -3.53629690529662e-15 walpha0 = -2.06600503969558e-16 palpha0 = 1.66574507412411e-21   alpha1 = 5.38602961623308e-10 lalpha1 = -3.53629690529662e-15 walpha1 = -2.06600503969558e-16 palpha1 = 1.66574507412411e-21   beta0 = -112.204824903227 lbeta0 = 0.000890239102227316 wbeta0 = 5.42663341730309e-05 pbeta0 = -4.1934018523918e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 3.26588221396565e-09 lagidl = -9.91886123424222e-15 wagidl = -9.85757084151413e-16 pagidl = 4.67220221727217e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.10455359771935 lkt1 = 1.76814845264831e-06 wkt1 = 2.72706865945636e-07 pkt1 = -8.32872537062056e-13   kt2 = -0.0355196086772416 wkt2 = -7.99094421033305e-9   at = -186853.8208675 wat = 0.0927264568598331   ute = -3.77471245901538 wute = 1.18477121016202e-6   ua1 = -2.55288928195512e-09 wua1 = 1.08190822841856e-15   ub1 = 1.14831103222126e-18 wub1 = -3.08047953753774e-25   uc1 = -1.63776641886191e-10 luc1 = 2.4046818956017e-16 wuc1 = 8.10059476359036e-17 puc1 = -1.13270665040439e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.101 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.924440585743439+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.25555270473803e-07 wvth0 = -6.12646108970582e-08 pvth0 = 3.84735263682512e-15   k1 = 0.566050075653426 lk1 = -4.83011508196845e-07 wk1 = -3.33736515584827e-08 pk1 = 1.64727307380771e-13   k2 = 0.0133550391597231 lk2 = 9.17154153153742e-08 wk2 = -2.63898482087518e-09 pk2 = -1.6361585557418e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -135636.656136208 lvsat = 0.93361800929343 wvsat = 0.0603734647755199 pvsat = -3.18403139849052e-7   ua = -1.46328288971607e-09 lua = 1.67139988104561e-15 wua = 2.41404724348221e-16 pua = -6.00140867399164e-22   ub = 1.36975361962089e-18 lub = -3.18514525684914e-24 wub = -2.67873665632178e-25 pub = 1.14123043743053e-30   uc = -1.70191068244708e-11 luc = -1.38647124805404e-16 wuc = -2.17831391986147e-17 puc = 4.72845204673094e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00282749503215887 lu0 = 5.7863088812259e-09 wu0 = 1.63528437165748e-09 pu0 = -1.24979965257867e-15   a0 = 1.21885073877942 la0 = -8.8142616280293e-08 wa0 = 1.65327236082022e-08 pa0 = 3.0060351769987e-14   keta = -0.0113884751456729 lketa = 9.58891493624642e-08 wketa = 7.3076541657624e-09 pketa = -3.27022464547034e-14   a1 = 0.0   a2 = 0.8   ags = 0.26392598028978 lags = -2.7358748852502e-08 wags = -1.32016413481672e-08 pags = 9.33048789790477e-15   b0 = -2.5321428544429e-07 lb0 = 1.07633854303033e-12 wb0 = 1.0239784293401e-13 pb0 = -4.95035483938513e-19   b1 = 2.23468957847141e-08 lb1 = -1.31823851157864e-13 wb1 = -8.79447698372983e-15 pb1 = 5.53741511259054e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.178923502316033+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.60862484894954e-07 wvoff = -1.03389650015954e-08 pvoff = -3.63317794308793e-14   nfactor = {-1.86496448053723+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.66685401672248e-05 wnfactor = 1.29508348016448e-06 pnfactor = -5.93425607842819e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.31170076923077e-05 wcit = -6.17866416080154e-12   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -3.06670429053246 lpclm = 1.18119724125614e-05 wpclm = 1.25491351001197e-06 ppclm = -4.02838105791926e-12   pdiblc1 = 0.39   pdiblc2 = 0.00322886884532153 lpdiblc2 = -1.21023268900568e-08 wpdiblc2 = -9.31124032898553e-10 ppdiblc2 = 4.12740418770412e-15   pdiblcb = -0.225   drout = 0.56   pscbe1 = 760363325.88905 lpscbe1 = 293.829194375776 wpscbe1 = 9.26833133988521 ppscbe1 = -0.000100208154874144   pscbe2 = 9.3750721445518e-09 lpscbe2 = 1.82534082957351e-15 wpscbe2 = 3.78081618274997e-17 ppscbe2 = -6.22518252267583e-22   pvag = 0.0   delta = 0.01   alpha0 = 3.89692469097189e-10 lalpha0 = -2.33568550965683e-15 walpha0 = -9.87973569843375e-17 palpha0 = 7.96567324721485e-22   alpha1 = 4.68014095746002e-10 lalpha1 = -2.96716443289736e-15 walpha1 = -1.25508336844227e-16 palpha1 = 1.01192828595707e-21   beta0 = -77.8427320716076 lbeta0 = 0.000613189986803572 wbeta0 = 2.81934132355265e-05 pbeta0 = -2.09123662117461e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.98506481106281e-09 lagidl = -3.18426461705364e-14 wagidl = -1.75318381055897e-15 pagidl = 1.08596861038213e-20   bgidl = -183651126.400764 lbgidl = 9543.35055046161 wbgidl = 403.674984180195 pbgidl = -0.00325468526710064   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.41947859399625 lkt1 = 4.30727469478032e-06 wkt1 = 3.57582832762902e-07 pkt1 = -1.51719673240969e-12   kt2 = -0.00352468221177527 lkt2 = -2.57963509927674e-07 wkt2 = -2.01705032278987e-08 pkt2 = 9.81993753582672e-14   at = -437790.979307098 lat = 2.02321546924712 wat = 0.185667467369573 pat = -7.49349723094226e-7   ute = -8.00430668315037 lute = 3.41016871160912e-05 wute = 2.74859306221923e-06 pute = -1.26085294896269e-11   ua1 = -6.60089653292633e-09 lua1 = 3.2637617085956e-14 wua1 = 2.68692322572467e-15 pua1 = -1.29406549078501e-20   ub1 = 2.67487905951955e-18 lub1 = -1.23081653864802e-23 wub1 = -9.9315114186668e-25 pub1 = 5.52373899840027e-30   uc1 = 1.01574348565114e-11 luc1 = -1.16189930708046e-15 wuc1 = 2.42376820559435e-17 puc1 = 3.44431310218639e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.102 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.815624689536858+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.16524324459113e-07 wvth0 = -8.14052918739652e-08 pvth0 = 8.56716485194886e-14   k1 = 0.435332593468791 lk1 = 4.80463021907745e-08 wk1 = 1.90375434337036e-08 pk1 = -4.82004050198966e-14   k2 = 0.0859180277667175 lk2 = -2.03081739592969e-07 wk2 = -2.6828192837735e-08 pk2 = 8.19104101217812e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 204216.23693826 lvsat = -0.44708126852084 wvsat = -0.0583411230648461 pvsat = 1.63891255865557e-7   ua = -2.12969462450208e-09 lua = 4.37878951843317e-15 wua = 4.45379277560614e-16 pua = -1.42881563831286e-21   ub = 1.17239861995464e-18 lub = -2.38336333571505e-24 wub = -1.65804284580323e-25 pub = 7.26559491332783e-31   uc = -6.10376402942689e-11 luc = 4.01842419732701e-17 wuc = -8.52754172869925e-18 puc = -6.56817352667283e-24   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.00118758543988802 lu0 = 2.20981273800215e-08 wu0 = 3.22205345951852e-09 pu0 = -7.69626804614829e-15   a0 = 1.49849164254337 la0 = -1.22422237826606e-06 wa0 = -7.61537504286554e-08 pa0 = 4.06611943278138e-13   keta = 0.0507840073616866 lketa = -1.5669514062627e-07 wketa = -1.11642047994409e-08 pketa = 4.23422297079722e-14   a1 = 0.0   a2 = 0.8   ags = -0.615618063429171 lags = 3.54591030583377e-06 wags = 2.36658146205628e-07 pags = -1.00575937969007e-12   b0 = -9.19136734464555e-08 lb0 = 4.2103254730467e-13 wb0 = 1.50930308134591e-14 pb0 = -1.40347636634704e-19   b1 = 1.21184747037519e-08 lb1 = -9.02694789943465e-14 wb1 = -5.58863785426785e-15 pb1 = 4.23499872566663e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.0605308842263133+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.2012386427583e-07 wvoff = -5.10797801042494e-08 pvoff = 1.29183404156136e-13   nfactor = {0.615622435760839+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.59081349876947e-06 wnfactor = 3.5997895234455e-07 pnfactor = -2.1352648897349e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.31170076923077e-05 wcit = -6.17866416080154e-12   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.1619898605 leta0 = -3.33095122881999e-7   etab = -0.1416766705 letab = 2.91196365286779e-7   dsub = 0.8693957 ldsub = -1.2569627278566e-6   voffl = 0.0   minv = 0.0   pclm = 0.165801325718038 lpclm = -1.32052773923126e-06 wpclm = 1.58409164980531e-07 ppclm = 4.26319161370583e-13   pdiblc1 = 0.39   pdiblc2 = 0.00287526665240015 lpdiblc2 = -1.0665769184211e-08 wpdiblc2 = -1.08327758272884e-09 ppdiblc2 = 4.74554898107951e-15   pdiblcb = -0.972376570248923 lpdiblcb = 3.03632045460294e-06 wpdiblcb = 2.54886949746147e-07 ppdiblcb = -1.03551340774279e-12   drout = 0.56   pscbe1 = 866399867.969509 lpscbe1 = -136.958890868891 wpscbe1 = -31.2771398880668 ppscbe1 = 6.4513417264443e-5   pscbe2 = 9.92226375164169e-09 lpscbe2 = -3.97700586670896e-16 wpscbe2 = -1.36691701344385e-16 ppscbe2 = 8.64115228493229e-23   pvag = 0.0   delta = 0.01   alpha0 = -3.90135392442842e-10 lalpha0 = 8.32472794094446e-16 walpha0 = 2.0232918260275e-16 palpha0 = -4.26800797813522e-22   alpha1 = -5.32894392303806e-10 lalpha1 = 1.09916442517634e-15 walpha1 = 2.51016025985133e-16 palpha1 = -5.1775389839928e-22   beta0 = 218.427839716425 lbeta0 = -0.000590450096424216 wbeta0 = -8.17017532942839e-05 pbeta0 = 2.37340617442875e-10   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -3.16108024617824e-09 lagidl = 5.31483029252324e-15 wagidl = 1.41370731683951e-15 pagidl = -2.00624613221059e-21   bgidl = 3367302252.80153 lbgidl = -4882.88758411404 wbgidl = -807.34996836039 pbgidl = 0.00166527072403894   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.129093081878613 lkt1 = -9.35094521398247e-07 wkt1 = -7.67795699068878e-08 pkt1 = 2.47460470447902e-13   kt2 = -0.0708597502728991 lkt2 = 1.55944963100339e-08 wkt2 = 5.30992517545232e-09 pkt2 = -5.31838132946583e-15   at = 173762.805276984 lat = -0.461306175047982 wat = -0.0411587092496908 pat = 1.72162921433905e-7   ute = 2.19730187460491 lute = -7.34375547177055e-06 wute = -9.14169168477292e-07 pute = 2.27194753376558e-12   ua1 = 2.86610796689899e-09 lua1 = -5.82339514120536e-15 wua1 = -9.87211264790143e-16 pua1 = 1.98602349042599e-21   ub1 = -7.01919742072287e-19 lub1 = 1.41054574322125e-24 wub1 = 4.84901941344051e-25 pub1 = -4.81055623468811e-31   uc1 = -6.14149379621297e-10 luc1 = 1.37443328107603e-15 wuc1 = 2.24396066866509e-16 puc1 = -4.68739749931389e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.103 pmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.03878304231691+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.43770574002425e-07 wvth0 = -2.28776569459063e-08 pvth0 = -3.5049675333255e-14   k1 = 0.319795735895534 lk1 = 2.86357015021961e-07 wk1 = 4.32784278952514e-08 pk1 = -9.82005744638945e-14   k2 = -0.0439928629055891 lk2 = 6.48774001215764e-08 wk2 = 2.19610743337677e-08 pk2 = -1.87241863383126e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -221235.289986053 lvsat = 0.430471218071272 wvsat = 0.0923994604835998 pvsat = -1.47031999903642e-7   ua = 2.95719609339844e-09 lua = -6.11362457815573e-15 wua = -1.08614317777817e-15 pua = 1.73016077592222e-21   ub = -2.10666071547509e-18 lub = 4.38014905379707e-24 wub = 8.01709135233483e-25 pub = -1.26907045388513e-30   uc = -1.13339951774826e-10 luc = 1.48064977120903e-16 wuc = 1.39156747617857e-18 puc = -2.70277050988037e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0207741687292226 lu0 = -2.32010213158444e-08 wu0 = -3.5894100065836e-09 pu0 = 6.35331533464566e-15   a0 = -0.250511714696515 la0 = 2.38333840850449e-06 wa0 = 6.35425795633532e-07 pa0 = -1.06111906845248e-12   keta = -0.0763066636061285 lketa = 1.05446906757443e-07 wketa = 3.04921357901756e-08 pketa = -4.35797213331132e-14   a1 = 0.0   a2 = 2.34014566561108 la2 = -3.1767629754247e-06 wa2 = -5.25254666120466e-07 pa2 = 1.08341023401739e-12   ags = 2.30827547412412 lags = -2.48502361267808e-06 wags = -7.58889917097594e-07 pags = 1.04769588650556e-12   b0 = 5.30847028255281e-08 lb0 = 1.21953386467778e-13 wb0 = -5.65003063151767e-14 pb0 = 7.32350107363148e-21   b1 = 7.72778067228481e-08 lb1 = -2.24669593271551e-13 wb1 = -3.60802707220142e-14 pb1 = 1.05243187891729e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.461792832405992+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.07534277993607e-07 wvoff = 9.39268317837359e-08 pvoff = -1.69912743775274e-13   nfactor = {-0.305145498588011+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.49002442933892e-06 wnfactor = 9.09250052180682e-07 pnfactor = -3.2682123325587e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.31170076923077e-05 wcit = -6.17866416080154e-12   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -0.519661301 leta0 = 1.07290446557204e-06 weta0 = 1.55096364853693e-23 peta0 = 6.66587464911755e-29   etab = -0.0556834575322843 letab = 1.13823496477477e-07 wetab = 1.08333774887346e-07 petab = -2.23453360766086e-13   dsub = 0.26   voffl = 0.0   minv = 0.0   pclm = -1.82807783656554 lpclm = 2.79212318830301e-06 wpclm = 8.13806585334293e-07 ppclm = -9.2552846295306e-13   pdiblc1 = 0.37861541905357 lpdiblc1 = 2.3482269274181e-08 wpdiblc1 = 5.10811475938829e-09 ppdiblc1 = -1.05361916110748e-14   pdiblc2 = -0.00519206926683768 lpdiblc2 = 5.97422444157386e-09 wpdiblc2 = 2.51113947439487e-09 ppdiblc2 = -2.66843222879202e-15   pdiblcb = 1.26975314049785 lpdiblcb = -1.58838148771235e-06 wpdiblcb = -5.09773899492294e-07 ppdiblcb = 5.41705117008693e-13   drout = -0.198321695714591 ldrout = 1.56414314580535e-06 wdrout = 1.92836719310074e-07 pdrout = -3.97752345044291e-13   pscbe1 = 738835324.266795 lpscbe1 = 126.160584424986 wpscbe1 = 29.41365725988 ppscbe1 = -6.06697271832045e-5   pscbe2 = 1.06057537027077e-08 lpscbe2 = -1.80749293235779e-15 wpscbe2 = -2.46965861025446e-16 ppscbe2 = 3.13867195025543e-22   pvag = 0.0   delta = 0.01   alpha0 = -7.84990915030732e-11 lalpha0 = 1.89679917596643e-16 walpha0 = -9.46893726815063e-18 palpha0 = 1.00620525607531e-23   alpha1 = -1.06267598376398e-10 lalpha1 = 2.19187788203498e-16 walpha1 = 1.29540664304629e-21 palpha1 = -1.37654832435342e-27   beta0 = -152.710909834686 lbeta0 = 0.000175074791672388 wbeta0 = 7.08814384721056e-05 pbeta0 = -7.73832720557671e-11   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 4.45969536991149e-10 lagidl = -2.1252076581337e-15 wagidl = -1.83452553225875e-16 pagidl = 1.28811650786134e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.571155007447362 lkt1 = -2.3280795366973e-08 wkt1 = 5.18410691953358e-08 pkt1 = -1.78373473486296e-14   kt2 = -0.0757114106170181 lkt2 = 2.56017152989067e-08 wkt2 = 9.6891208646387e-09 pkt2 = -1.43510767674179e-14   at = -216315.5972515 lat = 0.343284360986566 wat = 0.10425139777752 pat = -1.27765490904487e-7   ute = -4.14765666485134 lute = 5.74359712013641e-06 wute = 1.10600234135013e-06 pute = -1.89493498892184e-12   ua1 = -4.12748331666515e-09 lua1 = 8.60185199674281e-15 wua1 = 1.43344431134893e-15 pua1 = -3.00691268583036e-21   ub1 = 4.13100025016925e-18 lub1 = -8.55801868373586e-24 wub1 = -1.20075445993364e-24 pub1 = 2.9958433247498e-30   uc1 = 1.94800106319856e-10 luc1 = -2.94136668706654e-16 wuc1 = -4.56364766182228e-17 puc1 = 8.82396354968719e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.104 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.99939658343403+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.01917026108041e-07 wvth0 = -3.85143099597424e-08 pvth0 = -1.84335736479383e-14   k1 = 0.574912015551874 lk1 = 1.5260761840509e-08 wk1 = -6.97784658666406e-08 pk1 = 2.19379770094553e-14   k2 = -0.0261205274491204 lk2 = 4.58855773167855e-08 wk2 = 2.44191000893081e-08 pk2 = -2.13361779111286e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 334717.06290753 lvsat = -0.16030487830286 wvsat = -0.108248018033212 pvsat = 6.61836353725053e-8   ua = -1.45023313721359e-09 lua = -1.43012279539662e-15 wua = 2.27831690040424e-16 pua = 3.33881150333205e-22   ub = 6.28372411679186e-19 lub = 1.4737989216241e-24 wub = -1.17059829057066e-26 pub = -4.04704639575934e-31   uc = 4.31516589172005e-11 luc = -1.82289550816503e-17 wuc = -3.84613041679751e-17 puc = 1.53214707193966e-23   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.00114436600334333 lu0 = -2.34164700682154e-09 wu0 = 2.25606959736124e-09 pu0 = 1.41686579268928e-16   a0 = 3.35233854528087 la0 = -1.44518718605735e-06 wa0 = -9.41639829467647e-07 pa0 = 6.14730793273788e-13   keta = -0.0113011234102555 lketa = 3.63695495347806e-08 wketa = 1.07927635558483e-08 pketa = -2.26464198207722e-14   a1 = 0.0   a2 = -2.28029133122215 la2 = 1.73308895401617e-06 wa2 = 1.05050933224093e-06 pa2 = -5.91056469673374e-13   ags = 0.197825640476807 lags = -2.42379422350763e-07 wags = -8.27449349865456e-08 pags = 3.29198535005041e-13   b0 = 4.22424482975192e-07 lb0 = -2.70521098830901e-13 wb0 = -1.36351801380387e-13 pb0 = 9.21767340867368e-20   b1 = -2.49648667449949e-07 lb1 = 1.22734901390482e-13 wb1 = 1.21440669543137e-13 pb1 = -6.21445490297513e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.0656553538616086+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.29522077654237e-08 wvoff = -1.01969660037787e-07 pvoff = 3.82543125009648e-14   nfactor = {17.2524971380122+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.01673938267327e-05 wnfactor = -6.0560729973933e-06 pnfactor = 4.1334046221945e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 3.78772616402769e-05 lcit = -1.56848067347621e-11 wcit = -1.31313666530116e-11 pcit = 7.38820587091717e-18   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 0.109320535198286 letab = -6.15160163497523e-08 wetab = -2.1667189521375e-07 petab = 1.21910014498803e-13   dsub = 0.333447817503076 ldsub = -7.80484418958339e-08 wdsub = -5.45522942943789e-08 pdsub = 5.79693409043903e-14   voffl = 0.0   minv = 0.0   pclm = 1.06399395473597 lpclm = -2.81102195862045e-07 wpclm = -1.56652206294168e-07 ppclm = 1.05717926465424e-13   pdiblc1 = 1.08818968710778 lpdiblc1 = -7.30538311782403e-07 wpdiblc1 = -2.25629391294455e-07 ppdiblc1 = 2.34654250346969e-13   pdiblc2 = 0.00250126853213462 lpdiblc2 = -2.20100865045047e-09 wpdiblc2 = -1.24411138333461e-09 ppdiblc2 = 1.32204003216393e-15   pdiblcb = 0.365410157918769 lpdiblcb = -6.27392269390485e-07 wpdiblcb = -2.78108099688404e-07 ppdiblcb = 2.95528234836687e-13   drout = 1.83493315665746 ldrout = -5.96470724009573e-07 wdrout = -4.17787095391151e-07 pdrout = 2.51119724162189e-13   pscbe1 = 922329351.466411 lpscbe1 = -68.827141650358 wpscbe1 = -58.82731451976 ppscbe1 = 3.30984825867688e-5   pscbe2 = 4.22740139583817e-08 lpscbe2 = -3.54593896739268e-14 wpscbe2 = -1.14254805050777e-14 ppscbe2 = 1.21925816393519e-20   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 16.1233285347771 lbeta0 = -4.33488572006144e-06 wbeta0 = -4.46326727385587e-06 pbeta0 = 2.68087536870984e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -2.68344069420212e-09 lagidl = 1.20022257112105e-15 wagidl = 1.72059723834053e-15 pagidl = -7.35199154549205e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.687208025941646 lkt1 = 1.00041552099756e-07 wkt1 = 7.45018854779272e-08 pkt1 = -4.19175918415301e-14   kt2 = -0.0893541092237358 lkt2 = 4.0098965260952e-08 wkt2 = 2.23761123877231e-08 pkt2 = -2.78327560655252e-14   at = 114190.896063337 lat = -0.00792439805652689 wat = -0.0158367305867719 pat = -1.55282355712579e-10   ute = 2.62420964319068 lute = -1.45244534970875e-06 wute = -1.36789158582845e-06 pute = 7.33918706067357e-13   ua1 = 8.31988786513549e-09 lua1 = -4.62519762114345e-15 wua1 = -3.08031418410275e-15 pua1 = 1.78957861425943e-21   ub1 = -8.9161196037379e-18 lub1 = 5.30634666358034e-24 wub1 = 3.45994266194706e-24 pub1 = -1.95679054345126e-30   uc1 = -2.01636058974268e-10 luc1 = 1.27131465109164e-16 wuc1 = 7.94891625124736e-17 puc1 = -4.47236234176932e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.105 pmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.602265034183334+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.21524274499271e-07 wvth0 = -1.60412751900271e-07 pvth0 = 5.01511219285971e-14   k1 = 0.629285050676495 lk1 = -1.53315738959383e-08 wk1 = -6.92881578752786e-08 pk1 = 2.16621111018114e-14   k2 = 0.156069691937285 lk2 = -5.66215633383429e-08 wk2 = -3.03882571003219e-08 pk2 = 9.50052392333044e-15   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -68059.3591788521 lvsat = 0.066312442266978 wvsat = 0.0211167480093405 pvsat = -6.6018978641442e-9   ua = -7.01452097887e-09 lua = 1.70055698725726e-15 wua = 1.84827166701667e-15 pua = -5.77839957432759e-22   ub = 5.590382449893e-18 lub = -1.31801648225645e-24 wub = -1.64516348154414e-24 pub = 5.14340620542996e-31   uc = 2.41299109629358e-11 luc = -7.52659685615862e-18 wuc = -2.52732821402585e-17 puc = 7.90138838176614e-24   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = -0.0122256566561298 lu0 = 5.18083580225912e-09 wu0 = 5.64414826155623e-09 pu0 = -1.76457522419642e-15   a0 = 0.748277688809539 la0 = 1.99564061059633e-08 wa0 = 3.3971377160708e-07 pa0 = -1.06207434127694e-13   keta = 0.132511992490296 lketa = -4.45451743692739e-08 wketa = -6.6296003676947e-08 pketa = 2.07266499975534e-14   a1 = 0.0   a2 = 1.14549842976048 la2 = -1.94390545523577e-7   ags = -1.05178808414181 lags = 4.60700744441208e-07 wags = 1.13057236109632e-06 pags = -3.53459881828432e-13   b0 = -1.31396130314817e-07 lb0 = 4.10794233893639e-14 wb0 = 6.18401170467136e-14 pb0 = -1.93335705132504e-20   b1 = -7.09077022648896e-08 lb1 = 2.21684422206906e-14 wb1 = 2.47303456026418e-14 pb1 = -7.73164578851873e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {0.155598922667777+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.03557877431388e-07 wvoff = -7.64707723335012e-08 pvoff = 2.39076693208012e-14   nfactor = {-4.13902731691107+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.86829070953644e-06 wnfactor = 2.9041112923485e-06 pnfactor = -9.07935546217249e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 0.49   etab = 4.56432325650385e-05 letab = -3.38096839426685e-11 wetab = 8.69087811526264e-12 petab = -2.71709875219948e-18   dsub = -0.347099133666233 ldsub = 3.04853133616163e-07 wdsub = 1.09104588588758e-07 pdsub = -3.41102403672121e-14   voffl = 0.0   minv = 0.0   pclm = 0.473371630760217 lpclm = 5.12043672550275e-08 wpclm = 7.03177696819451e-08 ppclm = -2.1984006877824e-14   pdiblc1 = -1.05081865450095 lpdiblc1 = 4.72949063523649e-07 wpdiblc1 = 4.30826323551357e-07 ppdiblc1 = -1.34692680142449e-13   pdiblc2 = -0.0170152014278372 lpdiblc2 = 8.77969897488817e-09 wpdiblc2 = 2.48822276666922e-09 ppdiblc2 = -7.77912989325933e-16   pdiblcb = -1.40582031583754 lpdiblcb = 3.69169301902816e-07 wpdiblcb = 5.56216199376808e-07 ppdiblcb = -1.73894320140767e-13   drout = 1.20389181490977 ldrout = -2.41422885571342e-07 wdrout = 6.42273135420088e-08 pdrout = -2.00798988511466e-14   pscbe1 = 800088964.269279 lpscbe1 = -0.0500546785392544   pscbe2 = -5.82148656475319e-08 lpscbe2 = 2.10794725697853e-14 wpscbe2 = 2.30566885557441e-14 ppscbe2 = -7.20839699669072e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.32526294943312 lbeta0 = 6.15240304745327e-07 wbeta0 = 6.78686385128496e-07 pbeta0 = -2.12183154073802e-13   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.36338773673375e-09 lagidl = 4.57510615236967e-16 wagidl = 9.31496937744939e-16 pagidl = -2.91221339622702e-22   bgidl = 653150899.046399 lbgidl = 195.150484462332   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.506061026159999 lkt1 = -1.87863356338981e-9   kt2 = -0.018700497393889 lkt2 = 3.46558408230713e-10 wkt2 = -6.09724197756858e-08 pkt2 = 1.90622953738308e-14   at = 142063.218379028 lat = -0.0236064257395827 wat = -0.036262515118371 pat = 1.13370402015773e-8   ute = 0.32782863110708 lute = -1.60414129832055e-07 wute = -1.42836319999964e-07 pute = 4.46560614121489e-14   ua1 = -2.79847411997416e-10 lua1 = 2.13340235712048e-16 wua1 = 2.25907209376891e-16 pua1 = -7.06271781251724e-23   ub1 = 6.10203519889804e-19 lub1 = -5.35247260513088e-26 wub1 = -4.03812960747562e-26 pub1 = 1.26247276422196e-32   uc1 = 5.401768370832e-11 luc1 = -1.67090453662817e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.24e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.106 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.13223857783257+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 4.41655942401396e-8   k1 = -0.813567419469429 lk1 = 4.35758936665543e-7   k2 = 0.4650984288698 lk2 = -1.53235689595451e-07 wk2 = 2.64697796016969e-23 pk2 = 6.31088724176809e-30   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 232244.975086 lvsat = -0.0275741041889168   ua = 1.19798413021857e-09 lua = -8.66984185037974e-16   ub = -2.19204033057143e-19 lub = 4.98281016600118e-25   uc = -1.36281915230573e-14 luc = 2.15909380130795e-20   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0126037456797143 lu0 = -2.58177888521451e-09 wu0 = -3.30872245021211e-24   a0 = -0.881468577428572 la0 = 5.29477019290114e-7   keta = -0.253803388541297 lketa = 7.62316937256813e-08 wketa = -6.61744490042422e-24 pketa = 6.31088724176809e-30   a1 = 0.0   a2 = 0.0215210757579989 la2 = 1.5700748647705e-7   ags = -2.44893826583886 lags = 8.97502982946609e-7   b0 = 1.69201876171429e-07 lb0 = -5.28989361624831e-14   b1 = 2.22121223971429e-08 lb1 = -6.94435352199795e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.515090606662571+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.06125155639393e-7   nfactor = {4.14427546896857+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -7.21384506835397e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = 1.75980323404943 leta0 = -3.96988743486745e-7   etab = 0.342493169811143 letab = -1.07095919498416e-07 wetab = 2.1713491079517e-23 petab = -8.14745403673576e-30   dsub = 1.89976708939571 ldsub = -3.97602628629477e-7   voffl = 0.0   minv = 0.0   pclm = 0.675862949280857 lpclm = -1.21021135846287e-8   pdiblc1 = 1.47685958670628 lpdiblc1 = -3.172992064509e-7   pdiblc2 = 0.0377080596946343 lpdiblc2 = -8.32887193591908e-9   pdiblcb = -1.00488780626506 lpdiblcb = 2.43822563975097e-7   drout = -1.538265090594 ldrout = 6.15879565051547e-7   pscbe1 = 799682270.466856 lpscbe1 = 0.0770932584628099   pscbe2 = 3.76665057638886e-08 lpscbe2 = -8.8966876255384e-15   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 12.47154114788 lbeta0 = -9.93681818660703e-7   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = -1.55519579598486e-08 lagidl = 4.89339683265114e-15 wagidl = -1.97215226305253e-31 pagidl = 3.05628531213795e-37   bgidl = 2238746789.12 lbgidl = -300.567043418499   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.128944597999999 lkt1 = -1.19779559430476e-7   kt2 = 0.337380461485714 lkt2 = -1.10977880413971e-07 pkt2 = -3.15544362088405e-30   at = -32682.9420000003 lat = 0.031025864348996   ute = -0.369536229714286 lute = 5.76086255254149e-8   ua1 = 1.22407760542857e-09 lua1 = -2.56843873885977e-16   ub1 = 6.69020824e-19 lub1 = -7.19132503737119e-26   uc1 = -8.17431561011429e-11 luc1 = 2.57349520700691e-17 wuc1 = -2.31111593326468e-33 puc1 = -4.59177480789956e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8__model.107 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -3.1319e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 3.94789e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -5.722e-9   dwb = -1.7864e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -2.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25.0e+6   tnoib = .0e-6   epsrox = 3.9   toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.44996e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-2.08656567882462+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.75721613370646e-07 wvth0 = 5.94474098382219e-07 pvth0 = -1.44242006283265e-13   k1 = -4.37627881588999 lk1 = 1.30020810447024e-06 wk1 = 1.71766916823271e-06 pk1 = -4.16771811641649e-13   k2 = 1.26170387272372 lk2 = -3.46522441281278e-07 wk2 = -3.39111432012073e-07 pk2 = 8.22813196405455e-14   k3 = -15.845   dvt0 = 4.4955   dvt1 = 0.294   dvt2 = 0.015   dvt0w = -4.9772   dvt1w = 1147200.0   dvt2w = -0.00896   w0 = 0.0   k3b = 2.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 880276.084456222 lvsat = -0.184811076504289 wvsat = -0.273029062109399 pvsat = 6.62472255721004e-8   ua = 3.2076187616053e-09 lua = -1.35459791272839e-15 wua = -2.32886642805101e-15 pua = 5.65071492369441e-22   ub = -3.61906885549373e-18 lub = 1.32321741738649e-24 wub = 2.08934237271971e-24 pub = -5.06953854631966e-31   uc = 7.49533374653378e-13 luc = -1.63581058080838e-19 wuc = -5.93320302720995e-19 puc = 1.43962051611617e-25   rdsw = 547.88   prwb = -0.32348   prwg = 0.1376   wr = 1.0   u0 = 0.0191708116049653 lu0 = -4.17519862718557e-09 wu0 = -7.31609627784909e-09 pu0 = 1.77516296866475e-15   a0 = 10.1337238202022 la0 = -2.14322723368622e-06 wa0 = -1.97334093237014e-06 pa0 = 4.78807497148426e-13   keta = 1.35948240919999 lketa = -3.15212745666669e-07 wketa = -3.26912554478217e-07 pketa = 7.93214083934857e-14   a1 = 0.0   a2 = -5.05296529360328 la2 = 1.38827071016613e-06 wa2 = 2.25641580329822e-06 pa2 = -5.47492217680673e-13   ags = -14.8015178403205 lags = 3.89470818573969e-06 wags = 5.47424495760216e-06 pags = -1.32825984802267e-12   b0 = 1.31961705231629e-06 lb0 = -3.32033373671921e-13 wb0 = -2.93769881404763e-13 pb0 = 7.12797364842887e-20   b1 = 2.09018791404439e-07 lb1 = -5.22707500765902e-14 wb1 = -1.16944762240667e-13 pb1 = 2.83752432205509e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.686897998442072+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.47812157565988e-07 wvoff = 4.51963035607002e-07 pvoff = -1.09663407033612e-13   nfactor = {-21.3790224203458+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.47153744643208e-06 wnfactor = 8.82956297097534e-06 pnfactor = -2.14238750015151e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 0.00013   cdscb = 0.00078   cdscd = 0.0   eta0 = -2.18190401599902 leta0 = 5.59419220250509e-07 weta0 = 8.99142229271662e-07 peta0 = -2.18166072226018e-13   etab = -1.0931432955008 letab = 2.41244041171944e-07 wetab = 2.12650732829459e-07 petab = -5.15971485122744e-14   dsub = 0.268905946910668 ldsub = -1.89374273919029e-9   voffl = 0.0   minv = 0.0   pclm = 3.84670102149259 lpclm = -7.81467921749938e-07 wpclm = -1.48881647463989e-06 ppclm = 3.61243451773673e-13   pdiblc1 = 2.71344445084547 lpdiblc1 = -6.17341684715902e-07 wpdiblc1 = -1.22764103600396e-06 ppdiblc1 = 2.97872365693929e-13   pdiblc2 = 0.0620367624618421 lpdiblc2 = -1.42319397179488e-08 wpdiblc2 = -2.84728618432787e-08 ppdiblc2 = 6.90859825192945e-15   pdiblcb = 1.92341155235452 lpdiblcb = -4.66694135801643e-07 wpdiblcb = -6.55626368706527e-07 ppdiblcb = 1.59079870850214e-13   drout = -0.679330968135623 ldrout = 4.07469507446493e-07 wdrout = 7.91035753758735e-07 pdrout = -1.91935333220512e-13   pscbe1 = 744867507.64381 lpscbe1 = 13.3772376803227 wpscbe1 = 25.969730490945 ppscbe1 = -6.30124346686213e-6   pscbe2 = -8.28448691643609e-08 lpscbe2 = 2.03439513643022e-14 wpscbe2 = 1.14431698418282e-14 ppscbe2 = -2.77654784408152e-21   pvag = 0.0   delta = 0.01   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 30.7279174641248 lbeta0 = -5.4233724552817e-06 wbeta0 = -8.47196339336494e-06 pbeta0 = 2.05562025383929e-12   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 3.32635229634281e-08 lagidl = -6.95109382761086e-15 wagidl = -3.13778903634193e-15 pagidl = 7.61346856199933e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.114858387674985 lkt1 = -1.23197409331318e-07 wkt1 = -1.73161316498871e-07 pkt1 = 4.20155155126533e-14   kt2 = -0.12   at = 459360.135495277 lat = -0.0883624838883028 wat = -0.0495747623360452 pat = 1.20287211836933e-8   ute = -4.08285049135098 lute = 9.58599771340418e-07 wute = 1.41988776012302e-06 pute = -3.44518726340729e-13   ua1 = -1.20524261153093e-10 lua1 = 6.94076338176641e-17 wua1 = 1.82620811785608e-16 pua1 = -4.43107485300364e-23   ub1 = 3.7264e-19   uc1 = 2.70885236211404e-10 luc1 = -5.98260957838626e-17 wuc1 = -1.17157600884618e-16 puc1 = 2.8426885963442e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 1.5e+42   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 8.04e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0020386   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 6.5637e-11   cgso = 6.5637e-11   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 1.1939967e-11   cgdl = 1.1939967e-11   cf = 1.2e-11   clc = 1.0e-7   cle = 0.6   dlc = -2.0325e-8   dwc = 3.2175e-8   vfbcv = -0.14469   acde = 0.8   moin = 18.13   noff = 3.9   voffcv = -0.10701   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.000808127811   mjs = 0.34629   pbs = 0.6587   cjsws = 1.082848e-10   mjsws = 0.29781   pbsws = 0.7418   cjswgs = 2.6187824e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__pfet_01v8





















