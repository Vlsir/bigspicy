** Translated using xdm 2.6.0 on Nov_14_2022_16_05_05_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_01V8_LVT__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__nfet_01v8_lvt d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__nfet_01v8_lvt d g s b sky130_fd_pr__nfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__nfet_01v8_lvt__model.0 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4177611+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47213   k2 = -0.0324753   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 161140.0   ua = -1.3012667e-9   ub = 2.63804e-18   uc = 7.0152e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03165736   a0 = 1.9649815   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.503487   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11559919+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.1501979+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0047977   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.4345657e-5   alpha1 = 0.0   beta0 = 17.822982   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25364   kt2 = -0.034423   at = 333080.0   ute = -1.0777   ua1 = 2.6823e-9   ub1 = -2.4433e-18   uc1 = -1.9223e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.1 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.045100657e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = 1.060109905e-07 wvth0 = 9.147135941e-08 pvth0 = -7.317896269e-13   k1 = 5.492848205e-01 lk1 = -6.172543808e-07 wk1 = -5.325966398e-07 pk1 = 4.260882301e-12   k2 = -5.930836397e-02 lk2 = 2.146700126e-07 wk2 = 1.852275673e-07 pk2 = -1.481858510e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.325311799e+04 lvsat = 7.031130729e-01 wvsat = 6.066796310e-01 pvsat = -4.853561418e-6   ua = -1.339809067e-09 lua = 3.083468390e-16 wua = 2.660564193e-16 pua = -2.128505896e-21   ub = 2.668117703e-18 lub = -2.406277939e-25 wub = -2.076251841e-25 pub = 1.661044036e-30   uc = 6.984153296e-11 luc = 2.483800001e-18 wuc = 2.143141589e-18 puc = -1.714557205e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.125845003e-02 lu0 = 3.191361568e-09 wu0 = 2.753659594e-09 pu0 = -2.202984125e-14   a0 = 2.001829856e+00 la0 = -2.947944011e-07 wa0 = -2.543627269e-07 pa0 = 2.034953959e-12   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.913938252e-01 lags = 9.674787754e-08 wags = 8.347870195e-08 pags = -6.678467287e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.120495311e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.839799875e-08 wvoff = -2.450315329e-08 pvoff = 1.960302495e-13   nfactor = {1.254137926e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.315415186e-07 wnfactor = -7.174938444e-07 pnfactor = 5.740097842e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 3.413258877e-01 lpclm = -1.130636074e-06 wpclm = -9.755669500e-07 ppclm = 7.804735592e-12   pdiblc1 = 0.39   pdiblc2 = 2.875490026e-03 lpdiblc2 = 1.537807385e-08 wpdiblc2 = 1.326893856e-08 ppdiblc2 = -1.061542286e-13   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.386566658e-04 lalpha0 = -4.344992043e-10 walpha0 = -3.749067215e-10 palpha0 = 2.999330628e-15   alpha1 = 0.0   beta0 = 1.812552730e+01 lbeta0 = -2.420424426e-06 wbeta0 = -2.088458107e-06 pbeta0 = 1.670809299e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.532210306e-01 lkt1 = -3.351840832e-09 wkt1 = -2.892128788e-09 pkt1 = 2.313762319e-14   kt2 = -3.413616713e-02 lkt2 = -2.294721800e-09 wkt2 = -1.979995862e-09 pkt2 = 1.584037280e-14   at = 6.177481998e+05 lat = -2.277403956e+00 wat = -1.965053197e+00 pat = 1.572082841e-5   ute = -9.496457727e-01 lute = -1.024460070e-06 wute = -8.839532089e-07 pute = 7.071806882e-12   ua1 = 2.421249855e-09 lua1 = 2.088454672e-15 wua1 = 1.802018706e-15 pua1 = -1.441651906e-20   ub1 = -1.551862099e-18 lub1 = -7.131685954e-24 wub1 = -6.153560174e-24 pub1 = 4.922974287e-29   uc1 = -1.089195526e-11 luc1 = -6.665006577e-17 wuc1 = -5.750886858e-17 puc1 = 4.600827380e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.2 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.300877157e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.695147372e-09 wvth0 = -1.829427188e-07 pvth0 = 3.659229409e-13   k1 = 3.595646373e-01 lk1 = 1.416652445e-07 wk1 = 1.065193280e-06 pk1 = -2.130604924e-12   k2 = 6.261697871e-03 lk2 = -4.762367667e-08 wk2 = -3.704551346e-07 pk2 = 7.409862125e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.525746180e+05 lvsat = -8.142506882e-01 wvsat = -1.213359262e+00 pvsat = 2.426967263e-6   ua = -1.301518032e-09 lua = 1.551748471e-16 wua = -5.321128386e-16 pua = 1.064334760e-21   ub = 2.590971934e-18 lub = 6.797109765e-26 wub = 4.152503682e-25 pub = -8.305858627e-31   uc = 6.797964781e-11 luc = 9.931722285e-18 wuc = -4.286283177e-18 puc = 8.573445043e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.035081427e-02 lu0 = 6.822090648e-09 wu0 = -5.507319187e-09 pu0 = 1.101576738e-14   a0 = 1.913255540e+00 la0 = 5.952102035e-08 wa0 = 5.087254537e-07 pa0 = -1.017555196e-12   keta = 1.845489143e-01 lketa = -7.382334898e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.759922666e-01 lags = 3.566470059e-06 wags = -1.669574039e-07 pags = 3.339490341e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.224011073e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.301042801e-08 wvoff = 4.900630658e-08 pvoff = -9.802265944e-14   nfactor = {6.982521331e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.392115611e-06 wnfactor = 1.434987689e-06 pnfactor = -2.870269550e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081488e-01 leta0 = -3.180488942e-7   etab = -1.395071238e-01 letab = 2.780427440e-7   dsub = 8.370548752e-01 ldsub = -1.108276297e-6   voffl = 0.0   minv = 0.0   pclm = -1.127548607e-01 lpclm = 6.857800067e-07 wpclm = 1.951133900e-06 ppclm = -3.902667783e-12   pdiblc1 = 0.39   pdiblc2 = 4.747920834e-03 lpdiblc2 = 7.887966766e-09 wpdiblc2 = -2.653787713e-08 ppdiblc2 = 5.308119452e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.571458063e-05 lalpha0 = 3.830276776e-10 walpha0 = 7.498134429e-10 palpha0 = -1.499780598e-15   alpha1 = 0.0   beta0 = 1.374391235e+01 lbeta0 = 1.510693360e-05 wbeta0 = 4.176916215e-06 pbeta0 = -8.354688698e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.544879398e-01 lkt1 = 1.716055399e-09 wkt1 = 5.784257575e-09 pkt1 = -1.156970092e-14   kt2 = -3.976515447e-02 lkt2 = 2.022238152e-08 wkt2 = 3.959991724e-09 pkt2 = -7.920795247e-15   at = 4.547447476e+04 lat = 1.180826071e-02 wat = 3.930106394e+00 pat = -7.861018459e-6   ute = -1.242299076e+00 lute = 1.462131370e-07 wute = 1.767906418e-06 pute = -3.536175256e-12   ua1 = 2.634541885e-09 lua1 = 1.235242830e-15 wua1 = -3.604037412e-15 pua1 = 7.208813652e-21   ub1 = -2.902540144e-18 lub1 = -1.728696886e-24 wub1 = 1.230712035e-23 pub1 = -2.461676366e-29   uc1 = -2.035849816e-11 luc1 = -2.878195352e-17 wuc1 = 1.150177372e-16 puc1 = -2.300590530e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.3 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.291617716e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.547225364e-9   k1 = 4.289797110e-01 lk1 = 2.820867209e-9   k2 = -1.361539404e-02 lk2 = -7.865418038e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.853047423e+04 lvsat = 5.392657846e-2   ua = -9.429601312e-10 lua = -5.620144581e-16   ub = 2.563565418e-18 lub = 1.227897488e-25   uc = 5.933521056e-11 luc = 2.722236888e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.802997486e-02 lu0 = -8.537804747e-9   a0 = 2.198224308e+00 la0 = -5.104749335e-7   keta = -1.439316791e-01 lketa = -8.120496456e-8   a1 = 0.0   a2 = 0.38689047   ags = 7.351202806e-01 lags = 1.344017186e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.170973161e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.401758364e-9   nfactor = {1.002352380e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.838527771e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.500102500e-05 lcit = -1.000307521e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.934791593e-04 leta0 = -1.869774818e-10 weta0 = 8.271806126e-25   etab = -5.426287371e-04 letab = 8.526621309e-11 wetab = 8.271806126e-25   dsub = -5.984348308e-02 ldsub = 6.857042836e-7   voffl = 0.0   minv = 0.0   pclm = 2.292098176e-01 lpclm = 1.780547387e-9   pdiblc1 = 0.39   pdiblc2 = 6.973647912e-03 lpdiblc2 = 3.436056335e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.881059773e-04 lalpha0 = -1.246654715e-10   alpha1 = 0.0   beta0 = 2.119447407e+01 lbeta0 = 2.042828019e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.506093809e-01 lkt1 = -6.041857427e-9   kt2 = -4.635542289e-02 lkt2 = 3.340426936e-8   at = 3.048971878e+04 lat = 4.178084454e-2   ute = -1.328232595e+00 lute = 3.180977917e-7   ua1 = 3.274504592e-09 lua1 = -4.481377694e-17   ub1 = -3.911829725e-18 lub1 = 2.900891811e-25   uc1 = 1.241766698e-11 luc1 = -9.434100292e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.4 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.405433116e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.836647822e-9   k1 = 4.339008610e-01 lk1 = -2.101291677e-9   k2 = -1.525532726e-02 lk2 = -6.225148636e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.490951971e+04 lvsat = 5.754827527e-2   ua = -1.203528805e-09 lua = -3.013923677e-16   ub = 2.612519750e-18 lub = 7.382538090e-26   uc = 1.084869897e-10 luc = -2.193948633e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.324567759e-02 lu0 = -3.752526701e-9   a0 = 1.917502117e+00 la0 = -2.296951950e-7   keta = -4.409673090e-01 lketa = 2.158915577e-7   a1 = 0.0   a2 = 0.38689047   ags = 2.828531238e+00 lags = -7.498229206e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.149835578e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.875667690e-10   nfactor = {1.262960023e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.231917091e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.032425814e-04 leta0 = -3.967839054e-10   etab = -8.524558137e-04 letab = 3.951568042e-10   dsub = 2.512870653e-01 ldsub = 3.745099535e-7   voffl = 0.0   minv = 0.0   pclm = -5.514726820e-02 lpclm = 2.861959263e-7   pdiblc1 = 0.39   pdiblc2 = 1.029795449e-02 lpdiblc2 = 1.110682743e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.282973109e-05 lalpha0 = 9.631552873e-11   alpha1 = 0.0   beta0 = 1.841624069e+01 lbeta0 = 2.983085721e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.503774293e-01 lkt1 = -6.273856577e-9   kt2 = -7.439943100e-04 lkt2 = -1.221650956e-8   at = 7.236904387e+04 lat = -1.070658140e-4   ute = -1.004797786e+00 lute = -5.403321454e-9   ua1 = 4.070644646e-09 lua1 = -8.411170397e-16   ub1 = -4.740558503e-18 lub1 = 1.118987848e-24   uc1 = -1.724254986e-10 luc1 = 9.054005551e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.5 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.029766137e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.706609772e-8   k1 = 2.793768360e-01 lk1 = 7.519239825e-8   k2 = 2.293047540e-02 lk2 = -2.532587806e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.523796560e+04 lvsat = 2.737168499e-2   ua = -1.676308986e-09 lua = -6.490535728e-17   ub = 2.940894122e-18 lub = -9.042912150e-26   uc = 7.495628689e-11 luc = -5.167261156e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.179265608e-02 lu0 = -3.025718076e-9   a0 = 1.303272982e+00 la0 = 7.754528954e-8   keta = -1.408519794e-02 lketa = 2.362991351e-9   a1 = 0.0   a2 = 0.38689047   ags = 2.660090190e+00 lags = -6.655678660e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.190967010e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.344981570e-9   nfactor = {1.834614993e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.372470349e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -5.756722938e-03 leta0 = 2.884543647e-09 weta0 = 2.481541838e-24 peta0 = 9.737501799e-31   etab = 2.719813618e-02 letab = -1.363588956e-08 wetab = 1.271790192e-23 petab = -9.860761315e-31   dsub = 1.730440290e+00 ldsub = -3.653698854e-7   voffl = 0.0   minv = 0.0   pclm = 6.539922334e-01 lpclm = -6.851919806e-8   pdiblc1 = 0.39   pdiblc2 = 7.096194780e-03 lpdiblc2 = 1.712604490e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.545734797e-03 lalpha0 = 1.353283207e-09 walpha0 = 1.240770919e-24 palpha0 = 4.930380658e-31   alpha1 = 0.0   beta0 = 1.748592252e+01 lbeta0 = 3.448435521e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.529818574e-01 lkt1 = -4.971108619e-9   kt2 = -2.869288886e-02 lkt2 = 1.763667237e-9   at = 8.910788998e+04 lat = -8.479920332e-3   ute = -3.635657700e-01 lute = -3.261507820e-7   ua1 = 4.289527073e-09 lua1 = -9.506031243e-16   ub1 = -4.306647369e-18 lub1 = 9.019433299e-25   uc1 = 5.373579709e-11 luc1 = -2.258695540e-17 wuc1 = 2.465190329e-32 puc1 = -5.877471754e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.6 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.108344676e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.405267206e-8   k1 = 2.745297557e-01 lk1 = 7.640516197e-8   k2 = 2.103420774e-02 lk2 = -2.485142240e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.803744389e+05 lvsat = 1.066013683e-3   ua = -7.673197097e-10 lua = -2.923390192e-16   ub = 1.623316567e-18 lub = 2.392353704e-25   uc = 8.768374738e-11 luc = -8.351735406e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.645136350e-02 lu0 = -1.689299967e-9   a0 = 5.766152943e+00 la0 = -1.039089591e-6   keta = 2.854070882e-01 lketa = -7.257147609e-08 wketa = -2.646977960e-23 pketa = -4.417621069e-29   a1 = 0.0   a2 = 0.38689047   ags = -3.099011129e+00 lags = 7.753880794e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.723741828e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.567527388e-8   nfactor = {1.980480086e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.007508594e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.787339904e-01 leta0 = 4.616432086e-08 weta0 = -5.293955920e-23 peta0 = -6.310887242e-30   etab = -5.941179147e-02 letab = 8.034347384e-9   dsub = 1.369422259e-01 ldsub = 3.333129781e-8   voffl = 0.0   minv = 0.0   pclm = 9.769017293e-01 lpclm = -1.493127685e-7   pdiblc1 = -1.180357857e+00 lpdiblc1 = 3.929113876e-7   pdiblc2 = 1.454082521e-02 lpdiblc2 = -1.500792677e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.576463855e-03 lalpha0 = -1.429546506e-9   alpha1 = 0.0   beta0 = 3.711054217e+01 lbeta0 = -1.461742438e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.680736643e-01 lkt1 = -2.621556308e-8   kt2 = -3.720341457e-02 lkt2 = 3.893043323e-9   at = -8.429831643e+03 lat = 1.592450531e-2   ute = -1.057492229e+00 lute = -1.525269125e-7   ua1 = 1.705244192e-09 lua1 = -3.040026259e-16 wua1 = 1.577721810e-30   ub1 = -2.197171090e-18 lub1 = 3.741418174e-25   uc1 = -1.354486630e-10 luc1 = 2.474794243e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.7 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.635362363e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = 1.655270570e-8   k1 = 1.071428947e+00 lk1 = -6.720005673e-8   k2 = -2.099304360e-01 lk2 = 1.676956123e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.281421198e+05 lvsat = -7.541961255e-3   ua = -3.688485601e-09 lua = 2.340696803e-16   ub = 5.463068625e-18 lub = -4.527071491e-25   uc = 2.142995582e-10 luc = -3.116853759e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.953108929e-02 lu0 = -4.422319523e-10   a0 = 0.0   keta = 2.097403276e-01 lketa = -5.893594750e-8   a1 = 0.0   a2 = 0.38689047   ags = 9.669767833e-01 lags = 4.267672776e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.258881992e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.298267214e-9   nfactor = {5.438425398e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.478429588e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 6.574907252e-02 leta0 = 2.107250501e-9   etab = -8.906514992e-02 letab = 1.337803084e-8   dsub = 6.318557206e-01 ldsub = -5.585458851e-8   voffl = 0.0   minv = 0.0   pclm = 7.497989167e-02 lpclm = 1.321805627e-8   pdiblc1 = 4.081245638e+00 lpdiblc1 = -5.552558703e-7   pdiblc2 = 7.456255438e-02 lpdiblc2 = -1.096629497e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.888425476e-03 lalpha0 = -2.243285503e-10   alpha1 = 0.0   beta0 = 3.167255789e+01 lbeta0 = -4.817904819e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.915700017e-01 lkt1 = -3.960905600e-9   kt2 = 2.831994200e-02 lkt2 = -7.914593148e-9   at = 6.086296500e+04 lat = 3.437596887e-3   ute = -3.021925883e+00 lute = 2.014738543e-7   ua1 = -2.900311273e-09 lua1 = 5.259414967e-16 wua1 = 5.916456789e-31 pua1 = -2.115889831e-37   ub1 = 2.938405440e-18 lub1 = -5.513147512e-25 pub1 = -3.503246161e-46   uc1 = 5.856422250e-12 luc1 = -7.159404541e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.8 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.864309610e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.162706962e-7   k1 = 6.545513268e-01 wk1 = -1.259247122e-6   k2 = -9.591816850e-02 wk2 = 4.379435835e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -4.665572185e+04 wvsat = 1.434405556e+0   ua = -1.392394509e-09 wua = 6.290516222e-16   ub = 2.709154346e-18 wub = -4.908994837e-25   uc = 6.941794593e-11 wuc = 5.067145895e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.071419551e-02 wu0 = 6.510626727e-9   a0 = 2.052104066e+00 wa0 = -6.014035910e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.748944509e-01 wags = 1.973732226e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.072065390e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -5.793413429e-8   nfactor = {1.395948942e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.696409611e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 5.341444615e-01 wpclm = -2.306585852e-6   pdiblc1 = 0.39   pdiblc2 = 2.529147036e-04 wpdiblc2 = 3.137247111e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.127561208e-04 walpha0 = -8.864122953e-10   alpha1 = 0.0   beta0 = 1.853830626e+01 wbeta0 = -4.937854775e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.526494080e-01 wkt1 = -6.838016952e-9   kt2 = -3.374482548e-02 wkt2 = -4.681411606e-9   at = 1.006136464e+06 wat = -4.646081852e+0   ute = -7.749344451e-01 wute = -2.089978515e-6   ua1 = 2.065084985e-09 wua1 = 4.260610563e-15   ub1 = -3.356250215e-19 wub1 = -1.454919607e-23   uc1 = 4.745409231e-13 wuc1 = -1.359713371e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.9 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.864309610e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.162706962e-7   k1 = 6.545513268e-01 wk1 = -1.259247122e-6   k2 = -9.591816850e-02 wk2 = 4.379435835e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -4.665572185e+04 wvsat = 1.434405556e+0   ua = -1.392394509e-09 wua = 6.290516222e-16   ub = 2.709154346e-18 wub = -4.908994837e-25   uc = 6.941794593e-11 wuc = 5.067145895e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.071419551e-02 wu0 = 6.510626727e-9   a0 = 2.052104066e+00 wa0 = -6.014035910e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.748944509e-01 wags = 1.973732226e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.072065390e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -5.793413429e-8   nfactor = {1.395948942e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.696409611e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 5.341444615e-01 wpclm = -2.306585852e-6   pdiblc1 = 0.39   pdiblc2 = 2.529147036e-04 wpdiblc2 = 3.137247111e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.127561208e-04 walpha0 = -8.864122953e-10   alpha1 = 0.0   beta0 = 1.853830626e+01 wbeta0 = -4.937854775e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.526494080e-01 wkt1 = -6.838016952e-9   kt2 = -3.374482548e-02 wkt2 = -4.681411606e-9   at = 1.006136464e+06 wat = -4.646081852e+0   ute = -7.749344451e-01 wute = -2.089978515e-6   ua1 = 2.065084985e-09 wua1 = 4.260610563e-15   ub1 = -3.356250215e-19 wub1 = -1.454919607e-23   uc1 = 4.745409231e-13 wuc1 = -1.359713371e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.10 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.240709689e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.494527524e-07 wvth0 = 5.488866436e-07 pvth0 = -1.330531976e-12   k1 = 1.043597195e+00 lk1 = -1.556263229e-06 wk1 = -3.656656107e-06 pk1 = 9.590127411e-12   k2 = -2.364837733e-01 lk2 = 5.622912352e-07 wk2 = 1.305207143e-06 pk2 = -3.469232028e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.308736392e+05 lvsat = 3.368889343e-01 wvsat = 2.814160720e+00 pvsat = -5.519303506e-6   ua = -1.630478781e-09 lua = 9.523858948e-16 wua = 1.738690056e-15 pua = -4.438781213e-21   ub = 2.618246808e-18 lub = 3.636487852e-25 wub = 2.269730036e-25 pub = -2.871637113e-30   uc = 1.252660962e-10 luc = -2.234040501e-16 wuc = -3.997323452e-16 puc = 1.619280948e-21   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.405622741e-02 lu0 = 2.663323730e-08 wu0 = 3.794396215e-08 pu0 = -1.257397855e-13   a0 = 2.054922680e+00 la0 = -1.127503195e-08 wa0 = -4.691971468e-07 pa0 = -5.288528790e-13   keta = 1.046075667e-01 lketa = -4.184517114e-07 wketa = 5.518319249e-07 pketa = -2.207440825e-12   a1 = 0.0   a2 = 0.38689047   ags = -6.124457468e-01 lags = 4.349583696e-06 wags = 1.465271512e-06 pags = -5.071853076e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.696782395e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.095900904e-08 wvoff = -1.955882310e-07 pvoff = 5.506446057e-13   nfactor = {2.042699994e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.587136795e-06 wnfactor = -7.845682120e-06 pnfactor = 2.459835064e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.701199175e-06 lcit = 5.080740045e-11 wcit = 8.767586986e-11 pcit = -3.507214530e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081487e-01 leta0 = -3.180488942e-7   etab = -1.395071238e-01 letab = 2.780427440e-7   dsub = 1.188580884e+00 ldsub = -2.514452396e-06 wdsub = -2.426569980e-06 pdsub = 9.706777366e-12   voffl = 0.0   minv = 0.0   pclm = 3.789599667e-01 lpclm = 6.207697917e-07 wpclm = -1.443153885e-06 ppclm = -3.453904869e-12   pdiblc1 = 0.39   pdiblc2 = -7.953087507e-03 lpdiblc2 = 3.282569107e-08 wpdiblc2 = 6.113667541e-08 ppdiblc2 = -1.190629189e-13   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.081715920e-04 lalpha0 = -3.816814451e-10 walpha0 = -1.831107852e-09 palpha0 = 3.778975888e-15   alpha1 = 0.0   beta0 = 1.583256179e+01 lbeta0 = 1.082353257e-05 wbeta0 = -1.024094730e-05 pbeta0 = 2.121345723e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.795351465e-01 lkt1 = 1.075484655e-07 wkt1 = 1.786841237e-07 pkt1 = -7.421265945e-13   kt2 = -1.800341777e-02 lkt2 = -6.296885782e-08 wkt2 = -1.462604063e-07 pkt2 = 5.663450023e-13   at = 1.978398515e+06 lat = -3.889247516e+00 wat = -9.412790939e+00 pat = 1.906781352e-5   ute = -5.437118754e-01 lute = -9.249376793e-07 wute = -3.054413083e-06 pute = 3.857935983e-12   ua1 = -7.033509971e-10 lua1 = 1.107431146e-14 wua1 = 1.943730364e-14 pua1 = -6.070988351e-20   ub1 = 5.360017417e-18 lub1 = -2.278373736e-23 wub1 = -4.472898399e-23 pub1 = 1.207253385e-28   uc1 = 2.363201270e-11 luc1 = -9.263463439e-17 wuc1 = -1.886469997e-16 puc1 = 2.107134490e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.11 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.645061765e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.144645200e-08 wvth0 = -2.439810131e-07 pvth0 = 2.553658751e-13   k1 = 1.088850761e-01 lk1 = 3.133526258e-07 wk1 = 2.209600461e-06 pk1 = -2.143588308e-12   k2 = 1.032874557e-01 lk2 = -1.173208759e-07 wk2 = -8.069756955e-07 pk2 = 7.555666471e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.581588539e+03 lvsat = 6.195030038e-02 wvsat = 8.248267994e-02 pvsat = -5.538743150e-8   ua = -8.704844537e-10 lua = -5.677585588e-16 wua = -5.002967026e-16 pua = 3.965129746e-23   ub = 2.848812450e-18 lub = -9.752976448e-26 wub = -1.969048854e-24 pub = 1.520856788e-30   uc = -8.578631314e-11 luc = 1.987440344e-16 wuc = 1.001768073e-15 puc = -1.184007196e-21   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.397108366e-02 lu0 = -1.320055776e-08 wu0 = -4.101123646e-08 pu0 = 3.218679751e-14   a0 = 2.521661545e+00 la0 = -9.448484445e-07 wa0 = -2.232674316e-06 pa0 = 2.998462972e-12   keta = 1.582444314e-01 lketa = -5.257364364e-07 wketa = -2.085909604e-06 pketa = 3.068582969e-12   a1 = 0.0   a2 = 0.38689047   ags = 7.635827427e-01 lags = 1.597244631e-06 wags = -1.964752373e-07 pags = -1.748018920e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.423694708e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.985564197e-08 wvoff = 1.744526729e-07 pvoff = -1.895130603e-13   nfactor = {-3.405172368e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.179786227e-06 wnfactor = 9.269775248e-06 pnfactor = -9.636072768e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 4.040342335e-05 lcit = -3.541068105e-11 wcit = -1.753517397e-10 pcit = 1.753876868e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 7.612791964e-04 leta0 = -5.226119550e-10 weta0 = -1.158316944e-09 peta0 = 2.316871343e-15   etab = -5.907458106e-04 letab = 1.815102240e-10 wetab = 3.321502334e-10 petab = -6.643685577e-16   dsub = 1.879622467e-01 ldsub = -5.130099942e-07 wdsub = -1.710593040e-06 pdsub = 8.274676712e-12   voffl = 0.0   minv = 0.0   pclm = 1.255447267e+00 lpclm = -1.132384488e-06 wpclm = -7.084076063e-06 ppclm = 7.829095875e-12   pdiblc1 = 0.39   pdiblc2 = 1.061728113e-02 lpdiblc2 = -4.318853121e-09 wpdiblc2 = -2.515185433e-08 ppdiblc2 = 5.353182977e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.619443794e-04 lalpha0 = -8.919704317e-11 walpha0 = 1.805924639e-10 palpha0 = -2.448371418e-16   alpha1 = 0.0   beta0 = 2.067370522e+01 lbeta0 = 1.140253267e-06 wbeta0 = 3.594846489e-06 pbeta0 = -6.460966685e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.146162053e-01 lkt1 = -2.230272517e-08 wkt1 = -2.484594512e-07 pkt1 = 1.122481196e-13   kt2 = -1.436169478e-01 lkt2 = 1.882839531e-07 wkt2 = 6.713924162e-07 pkt2 = -1.069128261e-12   at = -5.287611467e+02 lat = 6.901271648e-02 wat = 2.141193262e-01 pat = -1.879805227e-7   ute = -1.415151130e+00 lute = 8.181194747e-07 wute = 5.999951699e-07 pute = -3.451629677e-12   ua1 = 3.761194344e-09 lua1 = 2.144305542e-15 wua1 = -3.359599890e-15 pua1 = -1.511140310e-20   ub1 = -4.724833787e-18 lub1 = -2.611967558e-24 wub1 = 5.612134523e-24 pub1 = 2.003278159e-29   uc1 = 1.732440977e-10 luc1 = -3.918894749e-16 wuc1 = -1.110178418e-15 puc1 = 2.053965200e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.12 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.362306525e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.165131587e-09 wvth0 = 2.977011277e-08 pvth0 = -1.844136971e-14   k1 = 4.509550580e-01 lk1 = -2.878748045e-08 wk1 = -1.177244395e-07 pk1 = 1.842136937e-13   k2 = -1.192256817e-02 lk2 = -2.087233952e-09 wk2 = -2.300590268e-08 pk2 = -2.856385954e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.674387031e+05 lvsat = -9.893978986e-02 wvsat = -1.052902852e+00 pvsat = 1.080230854e-6   ua = -5.975384403e-10 lua = -8.407605263e-16 wua = -4.183127249e-15 pua = 3.723236824e-21   ub = 2.190175441e-18 lub = 5.612422650e-25 wub = 2.915425870e-24 pub = -3.364619254e-30   uc = 1.388825644e-10 luc = -2.597090025e-17 wuc = -2.098194365e-16 puc = 2.782868901e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.925400679e-02 lu0 = -8.482513876e-09 wu0 = -4.147525610e-08 pu0 = 3.265091227e-14   a0 = 1.967143210e+00 la0 = -3.902164328e-07 wa0 = -3.426704785e-07 pa0 = 1.108071684e-12   keta = -7.017672566e-01 lketa = 3.344515540e-07 wketa = 1.800291606e-06 pketa = -8.184149121e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.457710894e-01 lags = 2.215182936e-06 wags = 1.851898600e-05 pags = -2.046731682e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.108344039e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.685889599e-09 wvoff = -2.864144353e-08 pvoff = 1.362269037e-14   nfactor = {9.862107925e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.527862186e-07 wnfactor = 1.910388870e-06 pnfactor = -2.275177716e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.422323427e-04 leta0 = -2.034996524e-10 weta0 = 2.492039543e-09 peta0 = -1.334233467e-15   etab = -7.578111693e-04 letab = 3.486098312e-10 wetab = -6.533281942e-10 petab = 3.213118930e-16   dsub = -1.650428431e+00 ldsub = 1.325757553e-06 wdsub = 1.312746600e-05 pdsub = -6.566424130e-12   voffl = 0.0   minv = 0.0   pclm = -6.068603868e-01 lpclm = 7.303049384e-07 wpclm = 3.808453589e-06 ppclm = -3.065666746e-12   pdiblc1 = 0.39   pdiblc2 = 4.724953150e-04 lpdiblc2 = 5.828012372e-09 wpdiblc2 = 6.782475167e-08 ppdiblc2 = -3.946383643e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.160757159e-04 lalpha0 = 1.888800462e-10 walpha0 = 5.746437034e-10 palpha0 = -6.389691618e-16   alpha1 = 0.0   beta0 = 1.812799754e+01 lbeta0 = 3.686482826e-06 wbeta0 = 1.989730935e-06 pbeta0 = -4.855522082e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.176063516e-01 lkt1 = -1.931196595e-08 wkt1 = -2.262174387e-07 pkt1 = 9.000154748e-14   kt2 = 9.092767469e-02 lkt2 = -4.630875111e-08 wkt2 = -6.328058642e-07 pkt2 = 2.353373797e-13   at = 9.160163287e+03 lat = 5.932180582e-02 wat = 4.363283743e-01 pat = -4.102351237e-7   ute = -2.523167320e-01 lute = -3.449533043e-07 wute = -5.194346617e-06 pute = 2.343899950e-12   ua1 = 9.461339951e-09 lua1 = -3.557008594e-15 wua1 = -3.721175406e-14 pua1 = 1.874769077e-20   ub1 = -1.229958909e-17 lub1 = 4.964340574e-24 wub1 = 5.217968581e-23 pub1 = -2.654431605e-29   uc1 = -5.338154579e-10 luc1 = 3.153150279e-16 wuc1 = 2.494660433e-15 puc1 = -1.551612643e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.13 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.235804563e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.685794020e-08 wvth0 = -1.422275015e-07 pvth0 = 6.759269692e-14   k1 = 2.609766475e-01 lk1 = 6.624067035e-08 wk1 = 1.270157651e-07 pk1 = 6.179341960e-14   k2 = 3.011652569e-02 lk2 = -2.311539889e-08 wk2 = -4.960501768e-08 pk2 = -1.525884923e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.803276194e+05 lvsat = 1.250351635e-01 wvsat = 2.454455011e+00 pvsat = -6.741670855e-7   ua = -1.879485214e-09 lua = -1.995243405e-16 wua = 1.402517372e-15 pua = 9.292694565e-22   ub = 3.105106033e-18 lub = 1.035894082e-25 wub = -1.133548259e-24 pub = -1.339302150e-30   uc = 1.392895125e-10 luc = -2.617445776e-17 wuc = -4.440896833e-16 puc = 1.450118378e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.958516011e-02 lu0 = -3.646108423e-09 wu0 = 1.523825641e-08 pu0 = 4.282529747e-15   a0 = 3.362407294e-01 la0 = 4.255691425e-07 wa0 = 6.675384959e-06 pa0 = -2.402394736e-12   keta = -1.398090560e-01 lketa = 5.335725228e-08 wketa = 8.678667629e-07 pketa = -3.520113434e-13   a1 = 0.0   a2 = 0.38689047   ags = 9.152393453e+00 lags = -2.289974604e-06 wags = -4.481610973e-05 pags = 1.121321474e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.240919189e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.945585679e-09 wvoff = 3.448178896e-08 pvoff = -1.795186614e-14   nfactor = {2.730206212e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.956901038e-08 wnfactor = -6.182230364e-06 pnfactor = 1.772790888e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.126486080e-02 leta0 = 5.652447413e-09 weta0 = 3.802246309e-08 peta0 = -1.910672898e-14   etab = -4.637919073e-02 letab = 2.316865199e-08 wetab = 5.079013445e-07 petab = -2.540602782e-13   dsub = 1.906712201e+00 ldsub = -4.535419765e-07 wdsub = -1.216797949e-06 pdsub = 6.086484180e-13   voffl = 0.0   minv = 0.0   pclm = 1.357918688e+00 lpclm = -2.524873787e-07 wpclm = -4.859176159e-06 ppclm = 1.269924993e-12   pdiblc1 = 0.39   pdiblc2 = 1.278350666e-02 lpdiblc2 = -3.300170571e-10 wpdiblc2 = -3.925928641e-08 ppdiblc2 = 1.410013484e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.932825733e-03 lalpha0 = 2.598242488e-09 walpha0 = 1.647799324e-08 palpha0 = -8.593904119e-15   alpha1 = 0.0   beta0 = 1.776203464e+01 lbeta0 = 3.869539297e-06 wbeta0 = -1.905990941e-06 pbeta0 = -2.906862521e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.704465940e-01 lkt1 = -4.290151247e-08 wkt1 = -5.697376216e-07 pkt1 = 2.618320606e-13   kt2 = 7.433412156e-03 lkt2 = -4.544503514e-09 wkt2 = -2.493784109e-07 pkt2 = 4.354505037e-14   at = 1.836829397e+05 lat = -2.797535955e-02 wat = -6.528477851e-01 pat = 1.345762371e-7   ute = 1.887776700e+00 lute = -1.415438739e-06 wute = -1.554092701e-05 pute = 7.519311198e-12   ua1 = 9.414788628e-09 lua1 = -3.533723390e-15 wua1 = -3.537947550e-14 pua1 = 1.783117587e-20   ub1 = -8.282970300e-18 lub1 = 2.955207769e-24 wub1 = 2.744839813e-23 pub1 = -1.417360230e-29   uc1 = 3.226412995e-10 luc1 = -1.130889244e-16 wuc1 = -1.856243927e-15 puc1 = 6.247314721e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.14 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.444500756e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -7.710012329e-08 wvth0 = -2.320471973e-07 pvth0 = 9.006603391e-14   k1 = 1.142270366e-01 lk1 = 1.029581568e-07 wk1 = 1.106563258e-06 pk1 = -1.832942609e-13   k2 = 4.065743768e-02 lk2 = -2.575278778e-08 wk2 = -1.354583714e-07 pk2 = 6.222089135e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.643995825e+05 lvsat = -1.125830608e-02 wvsat = -5.800222053e-01 pvsat = 8.507428633e-8   ua = -3.674750289e-09 lua = 2.496599578e-16 wua = 2.006987699e-14 pua = -3.741397258e-21   ub = 4.131589065e-18 lub = -1.532417787e-25 wub = -1.731450472e-23 pub = 2.709254061e-30   uc = -1.913226853e-11 luc = 1.346346398e-17 wuc = 7.373466852e-16 puc = -1.505894487e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.275696060e-03 lu0 = 4.075432094e-09 wu0 = 1.913987831e-07 pu0 = -3.979371483e-14   a0 = 7.281403632e+00 la0 = -1.312145341e-06 wa0 = -1.045971490e-05 pa0 = 1.884892923e-12   keta = 7.796836748e-01 lketa = -1.767044264e-07 wketa = -3.411971506e-06 pketa = 7.188255907e-13   a1 = 0.0   a2 = 0.38689047   ags = -3.176823019e+00 lags = 7.948570035e-07 wags = 5.371323683e-07 pags = -1.343932042e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.853131346e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.026343996e-08 wvoff = 8.931706720e-08 pvoff = -3.167192693e-14   nfactor = {1.686462216e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.415809561e-07 wnfactor = 2.029593591e-06 pnfactor = -2.818485244e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -9.822121506e-07 lcit = 1.496779391e-12 wcit = 4.129497119e-11 pcit = -1.033220827e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -7.044092267e-02 leta0 = 2.045859369e-08 weta0 = -7.475427150e-07 peta0 = 1.774456064e-13   etab = 1.892266051e-01 letab = -3.578109615e-08 wetab = -1.716340906e-06 petab = 3.024562541e-13   dsub = -5.182455423e-01 ldsub = 1.531945757e-07 wdsub = 4.522734956e-06 pdsub = -8.274114125e-13   voffl = 0.0   minv = 0.0   pclm = 7.922231862e-01 lpclm = -1.109475357e-07 wpclm = 1.274828595e-06 ppclm = -2.648336671e-13   pdiblc1 = -1.180367404e+00 lpdiblc1 = 3.929137763e-07 wpdiblc1 = 6.590027376e-11 ppdiblc1 = -1.648857800e-17   pdiblc2 = -1.766110476e-02 lpdiblc2 = 7.287376942e-09 wpdiblc2 = 2.222886345e-07 ppdiblc2 = -5.134046272e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.326699160e-02 lalpha0 = -4.457492808e-09 walpha0 = -1.014081254e-07 palpha0 = 2.090179220e-14   alpha1 = 0.0   beta0 = 5.320759326e+01 lbeta0 = -4.999116697e-06 wbeta0 = -1.111172998e-04 pbeta0 = 2.441835301e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.849129105e-01 lkt1 = 1.075903225e-08 wkt1 = 1.496832643e-06 pkt1 = -2.552341525e-13   kt2 = -1.002038800e-01 lkt2 = 2.238688516e-08 wkt2 = 4.348896926e-07 pkt2 = -1.276622505e-13   at = 7.137922269e+04 lat = 1.235919599e-04 wat = -5.509187097e-01 pat = 1.090730728e-7   ute = -6.511920208e+00 lute = 6.862074255e-07 wute = 3.765169817e-05 pute = -5.789749586e-12   ua1 = -1.511240728e-08 lua1 = 2.603103663e-15 wua1 = 1.160915754e-13 pua1 = -2.006763843e-20   ub1 = 1.260465879e-17 lub1 = -2.270981467e-24 wub1 = -1.021764396e-22 pub1 = 1.825918023e-29   uc1 = -4.794854885e-10 luc1 = 8.760720854e-17 wuc1 = 2.374872445e-15 puc1 = -4.339149996e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.15 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.261808222e-03+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.844520844e-08 wvth0 = 1.106367966e-06 pvth0 = -1.511230707e-13   k1 = 1.757160984e+00 lk1 = -1.931067552e-07 wk1 = -4.733580824e-06 pk1 = 8.691289035e-13   k2 = -3.858839874e-01 lk2 = 5.111210973e-08 wk2 = 1.214600327e-06 pk2 = -2.370652386e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.314291108e+05 lvsat = -2.333736221e-02 wvsat = -7.129859670e-01 pvsat = 1.090350210e-7   ua = -7.592208003e-09 lua = 9.556054250e-16 wua = 2.694723959e-14 pua = -4.980732384e-21   ub = 1.457224054e-17 lub = -2.034699378e-24 wub = -6.288024936e-23 pub = 1.092042907e-29   uc = 4.759058017e-10 luc = -7.574487147e-17 wuc = -1.805857435e-15 puc = 3.077086497e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.544602832e-02 lu0 = -4.344056247e-09 wu0 = -1.788897875e-07 pu0 = 2.693413703e-14   a0 = 0.0   keta = 7.448385221e-01 lketa = -1.704251557e-07 wketa = -3.693761433e-06 pketa = 7.696055444e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.157439939e+00 lags = 1.380114711e-08 wags = -1.314759546e-06 pags = 1.993269782e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-4.824761631e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.381370351e-08 wvoff = 2.461512451e-06 pvoff = -4.591533961e-13   nfactor = {-3.541774017e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.183735267e-06 wnfactor = 2.482413670e-05 pnfactor = -4.389539166e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.895849502e-05 lcit = -2.096635744e-12 wcit = -9.635493277e-11 pcit = 1.447299268e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -3.753414126e-01 leta0 = 7.540318648e-08 weta0 = 3.044829975e-06 peta0 = -5.059589142e-13   etab = -2.066582050e-01 letab = 3.555932605e-08 wetab = 8.117401554e-07 petab = -1.531165936e-13   dsub = 6.916945902e-01 ldsub = -6.484268592e-08 wdsub = -4.130653232e-07 pdsub = 6.204447687e-14   voffl = 0.0   minv = 0.0   pclm = 1.585903703e+00 lpclm = -2.539727333e-07 wpclm = -1.042984663e-05 ppclm = 1.844407333e-12   pdiblc1 = 1.047479473e+01 lpdiblc1 = -1.707404716e-06 wpdiblc1 = -4.413441362e-05 ppdiblc1 = 7.953237394e-12   pdiblc2 = 1.465488917e-01 lpdiblc2 = -2.230408546e-08 wpdiblc2 = -4.969188068e-07 ppdiblc2 = 7.826431424e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -7.599338496e-03 lalpha0 = 1.104774208e-09 walpha0 = 6.549365519e-08 palpha0 = -9.174743174e-15   alpha1 = 0.0   beta0 = 1.940732906e+01 lbeta0 = 1.091859912e-06 wbeta0 = 8.466638399e-05 pbeta0 = -1.086284573e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 1.678185793e-01 lkt1 = -8.884594587e-08 wkt1 = -3.171140999e-06 pkt1 = 5.859580376e-13   kt2 = 4.243726388e-01 lkt2 = -7.214442640e-08 wkt2 = -2.733935924e-06 pkt2 = 4.433759697e-13   at = -1.043488374e+05 lat = 3.179066703e-02 wat = 1.140450464e+00 pat = -1.957201091e-7   ute = -4.565978779e+00 lute = 3.355390502e-07 wute = 1.065853537e-05 pute = -9.254466846e-13   ua1 = -8.020861942e-09 lua1 = 1.325171735e-15 wua1 = 3.534695645e-14 pua1 = -5.517054365e-21   ub1 = 7.082001366e-18 lub1 = -1.275770986e-24 wub1 = -2.860307693e-23 pub1 = 5.000892409e-30   uc1 = -3.075770137e-10 luc1 = 5.662844184e-17 wuc1 = 2.163618471e-15 puc1 = -3.958459772e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.16 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4300959+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40031   k2 = -0.007497591   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 242950.0   ua = -1.26538932e-9   ub = 2.610042e-18   uc = 7.0441e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0320286876   a0 = 1.930681   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.514744   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05344474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.068446   pdiblc1 = 0.39   pdiblc2 = 0.006587   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.3789948e-5   alpha1 = 0.0   beta0 = 17.541356   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25403   kt2 = -0.03469   at = 68095.0   ute = -1.1969   ua1 = 2.9253e-9   ub1 = -3.2731e-18   uc1 = -2.6978e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.17 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4300959+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40031   k2 = -0.007497591   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 242950.0   ua = -1.26538932e-9   ub = 2.610042e-18   uc = 7.0441e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0320286876   a0 = 1.930681   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.514744   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05344474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.068446   pdiblc1 = 0.39   pdiblc2 = 0.006587   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.3789948e-5   alpha1 = 0.0   beta0 = 17.541356   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25403   kt2 = -0.03469   at = 68095.0   ute = -1.1969   ua1 = 2.9253e-9   ub1 = -3.2731e-18   uc1 = -2.6978e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.18 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.348908914e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.918094872e-8   k1 = 3.053202645e-01 lk1 = 3.799784147e-7   k2 = 2.703685742e-02 lk2 = -1.381448732e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.373039192e+05 lvsat = -7.774555195e-1   ua = -1.279438180e-09 lua = 5.619831946e-17   ub = 2.664072538e-18 lub = -2.161332265e-25   uc = 4.456034750e-11 luc = 1.035279155e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.171709326e-02 lu0 = 1.246441217e-9   a0 = 1.960192025e+00 la0 = -1.180501480e-7   keta = 2.160221400e-01 lketa = -8.641328445e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.166082049e-01 lags = 3.325579247e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.264569842e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.021584513e-8   nfactor = {4.586609309e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.379257167e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.500051250e-05 lcit = -2.000307511e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081487e-01 leta0 = -3.180488942e-7   etab = -1.395071237e-01 letab = 2.780427440e-7   dsub = 6.986576910e-01 ldsub = -5.546591887e-7   voffl = 0.0   minv = 0.0   pclm = 8.758796185e-02 lpclm = -7.657177150e-8   pdiblc1 = 0.39   pdiblc2 = 4.390374869e-03 lpdiblc2 = 8.786950832e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.152811310e-05 lalpha0 = 3.812917846e-10   alpha1 = 0.0   beta0 = 1.376491995e+01 lbeta0 = 1.510651835e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.434589166e-01 lkt1 = -4.228650077e-8   kt2 = -4.753331630e-02 lkt2 = 5.137589810e-8   at = 7.796101116e+04 lat = -3.946606718e-2   ute = -1.160396259e+00 lute = -1.460224483e-7   ua1 = 3.221030309e-09 lua1 = -1.182981862e-15   ub1 = -3.670740754e-18 lub1 = 1.590644532e-24   uc1 = -1.445571660e-11 luc1 = -5.009170068e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.19 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.152465392e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.011178289e-8   k1 = 5.550022385e-01 lk1 = -1.194367180e-7   k2 = -5.964050972e-02 lk2 = 3.522762991e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.323479792e+04 lvsat = 5.076760731e-2   ua = -9.714940930e-10 lua = -5.597529829e-16   ub = 2.451262530e-18 lub = 2.095304152e-25   uc = 1.164701301e-10 luc = -4.030639125e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.569093675e-02 lu0 = -6.702060391e-9   a0 = 2.070885784e+00 la0 = -3.394603591e-7   keta = -2.628996124e-01 lketa = 9.380883932e-8   a1 = 0.0   a2 = 0.38689047   ags = 7.239144964e-01 lags = 1.244320537e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.071475686e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.406944517e-9   nfactor = {1.531045475e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.342682403e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.274156191e-04 leta0 = -5.483685830e-11   etab = -5.236848544e-04 letab = 4.737456420e-11   dsub = -1.574055819e-01 ldsub = 1.157642850e-06 pdsub = 5.169878828e-26   voffl = 0.0   minv = 0.0   pclm = -1.748239372e-01 lpclm = 4.483058211e-07 wpclm = 6.776263578e-21 ppclm = -6.462348536e-27   pdiblc1 = 0.39   pdiblc2 = 5.539135062e-03 lpdiblc2 = 6.489194950e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.984059022e-04 lalpha0 = -1.386295324e-10   alpha1 = 0.0   beta0 = 2.139950283e+01 lbeta0 = -1.642124833e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.647800369e-01 lkt1 = 3.601107076e-10   kt2 = -8.063174690e-03 lkt2 = -2.757247651e-8   at = 4.270181738e+04 lat = 3.105954853e-2   ute = -1.294012423e+00 lute = 1.212372715e-7   ua1 = 3.082892906e-09 lua1 = -9.066787370e-16   ub1 = -3.591746800e-18 lub1 = 1.432640432e-24   uc1 = -5.090033679e-11 luc1 = 2.280501086e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.20 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.422412225e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.888434362e-9   k1 = 4.271865560e-01 lk1 = 8.405166706e-9   k2 = -1.656744773e-02 lk2 = -7.854262062e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -4.514182485e+04 lvsat = 1.191582473e-1   ua = -1.442109616e-09 lua = -8.904098402e-17   ub = 2.778798380e-18 lub = -1.180725799e-25   uc = 9.652013131e-11 luc = -2.035230268e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.088017455e-02 lu0 = -1.890311986e-9   a0 = 1.897958222e+00 la0 = -1.664973469e-7   keta = -3.382893351e-01 lketa = 1.692140169e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.884744551e+00 lags = -1.917157488e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.166170962e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.064524369e-9   nfactor = {1.371917293e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.934290432e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 9.453738564e-04 leta0 = -4.728806826e-10   etab = -8.897177856e-04 letab = 4.134825322e-10   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 1.620643752e-01 lpclm = 1.113484466e-7   pdiblc1 = 0.39   pdiblc2 = 1.416627674e-02 lpdiblc2 = -2.139715296e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.545663987e-08 lalpha0 = 5.987251099e-11   alpha1 = 0.0   beta0 = 1.852972316e+01 lbeta0 = 2.706155490e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.632795326e-01 lkt1 = -1.140701196e-9   kt2 = -3.683549405e-02 lkt2 = 1.205741176e-9   at = 9.725463090e+04 lat = -2.350444832e-2   ute = -1.301052562e+00 lute = 1.282788538e-7   ua1 = 1.948306520e-09 lua1 = 2.281402392e-16   ub1 = -1.764538173e-18 lub1 = -3.949427737e-25   uc1 = -3.014483804e-11 luc1 = 2.045257232e-18 wuc1 = -3.155443621e-30   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.21 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.794598356e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.003441156e-07 wvth0 = 2.312630217e-06 pvth0 = -1.156789198e-12   k1 = 2.866210632e-01 lk1 = 7.871672903e-8   k2 = -1.067414665e-03 lk2 = -1.560745610e-08 wk2 = 1.048477915e-07 pk2 = -5.244538956e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.928928776e+04 lvsat = 1.112287290e-01 wvsat = 1.211072196e+00 pvsat = -6.057843676e-7   ua = -1.212306653e-08 lua = 5.253627070e-15 wua = 5.213856589e-14 pua = -2.607997135e-20   ub = 7.973614508e-18 lub = -2.716545581e-24 wub = -2.524707599e-23 pub = 1.262871365e-29   uc = 4.962804075e-11 luc = 3.103355479e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -9.435052538e-02 lu0 = 6.075071027e-08 wu0 = 6.290867492e-07 pu0 = -3.146723374e-13   a0 = 1.683997416e+00 la0 = -5.947308197e-8   keta = 3.541278369e-02 lketa = -1.771365147e-8   a1 = 0.0   a2 = 0.38689047   ags = 1.040446408e-01 lags = -2.603248936e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.171300640e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.321113416e-9   nfactor = {-4.887243417e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.524292526e-06 wnfactor = 3.154669295e-05 pnfactor = -1.577981355e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -3.588146411e-03 leta0 = 1.794808955e-9   etab = 5.616582166e-02 letab = -2.812598357e-08 wetab = -1.164670302e-21 petab = 5.585135209e-28   dsub = 1.661041340e+00 ldsub = -3.306561834e-7   voffl = 0.0   minv = 0.0   pclm = 3.768535958e-01 lpclm = 3.909804463e-9   pdiblc1 = 0.39   pdiblc2 = 4.857077532e-03 lpdiblc2 = 2.516792696e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.605927627e-03 lalpha0 = 8.631377997e-10 walpha0 = 5.293955920e-23 palpha0 = 1.262177448e-29   alpha1 = 0.0   beta0 = 1.737721608e+01 lbeta0 = 3.282645294e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.854763180e-01 lkt1 = 9.962241845e-9   kt2 = -4.291595688e-02 lkt2 = 4.247219086e-9   at = 5.187331774e+04 lat = -8.044885751e-4   ute = -1.249928231e+00 lute = 1.027062079e-7   ua1 = 2.271691268e-09 lua1 = 6.638157129e-17   ub1 = -2.741153258e-18 lub1 = 9.356497492e-26   uc1 = -5.213336592e-11 luc1 = 1.304402882e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.22 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.265167068e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.594197858e-07 wvth0 = -8.259393631e-06 pvth0 = 1.488384029e-12   k1 = 3.376415721e-01 lk1 = 6.595114259e-8   k2 = 8.891101270e-02 lk2 = -3.812050852e-08 wk2 = -3.744563983e-07 pk2 = 6.747891526e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.020560673e+06 lvsat = -1.514489805e-01 wvsat = -4.325257841e+00 pvsat = 7.794330893e-7   ua = 3.797287878e-08 lua = -7.280628928e-15 wua = -1.862091639e-13 pua = 3.355582238e-20   ub = -1.756909765e-17 lub = 3.674368714e-24 wub = 9.016812855e-23 pub = -1.624874761e-29   uc = 1.297376366e-10 luc = -1.694046594e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.909829075e-01 lu0 = -8.570264130e-08 wu0 = -2.246738390e-06 pu0 = 4.048734916e-13   a0 = 5.169592736e+00 la0 = -9.315864589e-7   keta = 9.080843526e-02 lketa = -3.157392047e-8   a1 = 0.0   a2 = 0.38689047   ags = -3.068376279e+00 lags = 7.677230868e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.672800661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.386889470e-8   nfactor = {2.484359535e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.914511988e-06 wnfactor = -1.126667606e-04 pnfactor = 2.030311359e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 7.355220655e-06 lcit = -5.892879839e-13   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.213694008e-01 leta0 = 5.628476762e-08 peta0 = 1.211690350e-27   etab = -1.573017145e-01 letab = 2.528466131e-8   dsub = 3.948922493e-01 ldsub = -1.385935017e-8   voffl = 0.0   minv = 0.0   pclm = 1.049610404e+00 lpclm = -1.644173128e-7   pdiblc1 = -1.180354099e+00 lpdiblc1 = 3.929104472e-7   pdiblc2 = 2.721885279e-02 lpdiblc2 = -3.078235281e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.792744805e-03 lalpha0 = -2.374320360e-10   alpha1 = 0.0   beta0 = 3.077306930e+01 lbeta0 = -6.906416019e-8   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -8.270319286e-02 lkt1 = -4.077260793e-8   kt2 = -1.239988143e-02 lkt2 = -3.388055572e-9   at = -3.985097293e+04 lat = 2.214538757e-2   ute = 1.089937704e+00 lute = -4.827399485e-7   ua1 = 8.326420291e-09 lua1 = -1.448541904e-15   ub1 = -8.024710231e-18 lub1 = 1.415537347e-24   uc1 = 0.0   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.23 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-6.551381494e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.668338159e-07 wvth0 = 4.367396620e-06 pvth0 = -7.870267080e-13   k1 = 8.014535233e-01 lk1 = -1.763009007e-8   k2 = -3.959591819e-01 lk2 = 4.925552489e-08 wk2 = 1.264502362e-06 pk2 = -2.278696482e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 9.910372895e+04 lvsat = 1.460216812e-02 wvsat = 4.377123562e-01 pvsat = -7.887795514e-8   ua = -7.637128700e-09 lua = 9.385224709e-16 wua = 2.716973001e-14 pua = -4.896121196e-21   ub = -5.664487347e-18 lub = 1.529098415e-24 wub = 3.735145439e-23 pub = -6.730918839e-30   uc = 1.113041423e-10 luc = -1.361865811e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -4.300870820e-02 lu0 = 1.052531781e-08 wu0 = 2.592229843e-07 pu0 = -4.671327788e-14   a0 = 0.0   keta = -9.299542930e-04 lketa = -1.504220398e-8   a1 = 0.0   a2 = 0.38689047   ags = 8.919906833e-01 lags = 5.404515841e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {1.450189676e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.888912392e-8   nfactor = {-7.723165518e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.447995853e-05 wnfactor = 3.898071705e-04 pnfactor = -7.024520116e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.955148609e-07 lcit = 8.254538097e-13   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.394081463e-01 leta0 = -2.674965025e-8   etab = -4.276829766e-02 letab = 4.645166929e-9   dsub = 6.082969202e-01 ldsub = -5.231593890e-8   voffl = 0.0   minv = 0.0   pclm = -5.198768067e-01 lpclm = 1.184121300e-7   pdiblc1 = 1.564079999e+00 lpdiblc1 = -1.016502994e-7   pdiblc2 = 4.622124783e-02 lpdiblc2 = -6.502561881e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 5.623795789e-03 lalpha0 = -7.476015785e-10   alpha1 = 0.0   beta0 = 3.650142714e+01 lbeta0 = -1.101342885e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.724331083e-01 lkt1 = 2.945867149e-8   kt2 = -1.276075758e-01 lkt2 = 1.737294700e-8   at = 1.259075070e+05 lat = -7.725119304e-3   ute = -2.414026133e+00 lute = 1.486918549e-7   ua1 = -8.843301617e-10 lua1 = 2.112813814e-16   ub1 = 1.307055287e-18 lub1 = -2.660934577e-25   uc1 = 1.292564093e-10 luc1 = -2.329265124e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.24 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.359699790e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.880037431e-8   k1 = 2.484262163e-01 wk1 = 7.446801162e-7   k2 = 5.252807771e-02 wk2 = -2.943034527e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.500415345e+05 wvsat = -5.250655099e-1   ua = -1.506612665e-09 wua = 1.182708410e-15   ub = 2.908071475e-18 wub = -1.461226597e-24   uc = 7.253527625e-11 wuc = -1.026815269e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.213053522e-02 wu0 = -4.993548116e-10   a0 = 2.287114591e+00 wa0 = -1.747579642e-6   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.021348355e-01 wags = 6.182222939e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.249036685e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 2.941902722e-8   nfactor = {5.330374098e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.551536324e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.731899497e-05 wcit = -3.588473960e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.241226130e-01 wpclm = 9.441562067e-7   pdiblc1 = 0.39   pdiblc2 = 6.404757025e-03 wpdiblc2 = 8.935300161e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.642123509e-05 walpha0 = 3.612850464e-11   alpha1 = 0.0   beta0 = 1.716897432e+01 wbeta0 = 1.825772489e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.514390758e-01 wkt1 = -1.270319782e-8   kt2 = -3.455825809e-02 wkt2 = -6.459253128e-10   at = -2.984183114e+05 wat = 1.797000105e+0   ute = -1.103070484e+00 wute = -4.600423617e-7   ua1 = 4.155476675e-09 wua1 = -6.031507032e-15   ub1 = -5.006823530e-18 wub1 = 8.500377117e-24   uc1 = 2.069627256e-12 wuc1 = -1.424193545e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.25 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.359699790e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.880037431e-8   k1 = 2.484262163e-01 wk1 = 7.446801162e-7   k2 = 5.252807771e-02 wk2 = -2.943034527e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.500415345e+05 wvsat = -5.250655099e-1   ua = -1.506612665e-09 wua = 1.182708410e-15   ub = 2.908071475e-18 wub = -1.461226597e-24   uc = 7.253527625e-11 wuc = -1.026815269e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.213053522e-02 wu0 = -4.993548116e-10   a0 = 2.287114591e+00 wa0 = -1.747579642e-6   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.021348355e-01 wags = 6.182222939e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.249036685e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 2.941902722e-8   nfactor = {5.330374098e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.551536324e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.731899497e-05 wcit = -3.588473960e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.241226130e-01 wpclm = 9.441562067e-7   pdiblc1 = 0.39   pdiblc2 = 6.404757025e-03 wpdiblc2 = 8.935300161e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.642123509e-05 walpha0 = 3.612850464e-11   alpha1 = 0.0   beta0 = 1.716897432e+01 wbeta0 = 1.825772489e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.514390758e-01 wkt1 = -1.270319782e-8   kt2 = -3.455825809e-02 wkt2 = -6.459253128e-10   at = -2.984183114e+05 wat = 1.797000105e+0   ute = -1.103070484e+00 wute = -4.600423617e-7   ua1 = 4.155476675e-09 wua1 = -6.031507032e-15   ub1 = -5.006823530e-18 wub1 = 8.500377117e-24   uc1 = 2.069627256e-12 wuc1 = -1.424193545e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.26 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.608289775e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.944109022e-08 wvth0 = -1.271733985e-07 pvth0 = 3.935122634e-13   k1 = -7.577401948e-02 lk1 = 1.296867404e-06 wk1 = 1.868490031e-06 pk1 = -4.495470039e-12   k2 = 1.804586243e-01 lk2 = -5.117484123e-07 wk2 = -7.522207863e-07 pk2 = 1.831763208e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.361221084e+05 lvsat = -1.144380942e+00 wvsat = -9.747976285e-01 pvsat = 1.799020670e-6   ua = -1.736878994e-09 lua = 9.211125222e-16 wua = 2.242814015e-15 pua = -4.240639739e-21   ub = 3.246288191e-18 lub = -1.352936198e-24 wub = -2.854580062e-24 pub = 5.573699498e-30   uc = 3.790710812e-11 luc = 1.385197713e-16 wuc = 3.262056656e-17 puc = -1.715636692e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.100852886e-02 lu0 = 4.488255464e-09 wu0 = 3.474062946e-09 pu0 = -1.589448558e-14   a0 = 2.531836372e+00 la0 = -9.789372890e-07 wa0 = -2.802749368e-06 pa0 = 4.220895217e-12   keta = 1.635981251e-01 lketa = -6.544260379e-07 wketa = 2.570328482e-07 pketa = -1.028184085e-12   a1 = 0.0   a2 = 0.38689047   ags = 2.019838575e-01 lags = 1.200665443e-06 wags = -2.542636138e-06 pags = 1.041836738e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.480502762e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.259117589e-08 wvoff = 1.058710470e-07 pvoff = -3.058237517e-13   nfactor = {-1.022661172e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.223113245e-06 wnfactor = 7.262863017e-06 pnfactor = -1.884627259e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.963925265e-05 lcit = -4.928355634e-11 wcit = -7.177315739e-11 pcit = 1.435610283e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081488e-01 leta0 = -3.180488942e-7   etab = -1.394956610e-01 letab = 2.779968907e-07 wetab = -5.620126226e-11 petab = 2.248165703e-16   dsub = 5.857477084e-01 ldsub = -1.029961120e-07 wdsub = 5.535931280e-07 pdsub = -2.214485998e-12   voffl = 0.0   minv = 0.0   pclm = -1.007351989e-01 lpclm = -9.355445062e-08 wpclm = 9.233409244e-07 ppclm = 8.326539640e-14   pdiblc1 = 0.39   pdiblc2 = 2.854271827e-03 lpdiblc2 = 1.420266864e-08 wpdiblc2 = 7.531451770e-09 ppdiblc2 = -2.655304779e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.736173475e-05 lalpha0 = 3.351490549e-10 walpha0 = -2.042758640e-11 palpha0 = 2.262359582e-16   alpha1 = 0.0   beta0 = 1.324252449e+01 lbeta0 = 1.570660424e-05 wbeta0 = 2.561284079e-06 pbeta0 = -2.942197138e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.219684103e-01 lkt1 = -1.178887033e-07 wkt1 = -1.053670925e-07 pkt1 = 3.706745750e-13   kt2 = -6.834775718e-02 lkt2 = 1.351649232e-07 wkt2 = 1.020523710e-07 pkt2 = -4.108142385e-13   at = -6.777987810e+05 lat = 1.517599652e+00 wat = 3.705460031e+00 pat = -7.634230937e-6   ute = -9.389103874e-01 lute = -6.566740410e-07 wute = -1.085936368e-06 pute = 2.503704333e-12   ua1 = 5.094466190e-09 lua1 = -3.756150553e-15 wua1 = -9.185381187e-15 pua1 = 1.261614316e-20   ub1 = -6.588213473e-18 lub1 = 6.325883958e-24 wub1 = 1.430425204e-23 pub1 = -2.321668949e-29   uc1 = 2.316626015e-11 luc1 = -8.439085640e-17 wuc1 = -1.844590471e-16 puc1 = 1.681673885e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.27 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.891043541e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.402286013e-08 wvth0 = 1.281740877e-07 pvth0 = -1.172350553e-13   k1 = 7.127430665e-01 lk1 = -2.803284139e-07 wk1 = -7.733969702e-07 pk1 = 7.888455495e-13   k2 = -1.251850465e-01 lk2 = 9.960158642e-08 wk2 = 3.213622422e-07 pk2 = -3.156229338e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.006984299e+04 lvsat = 7.841679403e-03 wvsat = -1.806007526e-01 pvsat = 2.104641075e-7   ua = -9.568824803e-10 lua = -6.390404048e-16 wua = -7.164015246e-17 pua = 3.887430581e-22   ub = 2.255323699e-18 lub = 6.291959338e-25 wub = 9.606802488e-25 pub = -2.057603251e-30   uc = 1.342757448e-10 luc = -5.423725761e-17 wuc = -8.730021641e-17 puc = 6.830248051e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.498453278e-02 lu0 = -3.464567463e-09 wu0 = 3.463470404e-09 pu0 = -1.587329832e-14   a0 = 2.021442021e+00 la0 = 4.195604340e-08 wa0 = 2.424207924e-07 pa0 = -1.870069365e-12   keta = -1.819749615e-01 lketa = 3.679097766e-08 wketa = -3.967703268e-07 pketa = 2.795562950e-13   a1 = 0.0   a2 = 0.38689047   ags = -2.952329577e-01 lags = 2.195201003e-06 wags = 4.996839201e-06 pags = -4.662128887e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.876460842e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.599231317e-08 wvoff = -9.013091822e-08 pvoff = 8.622035909e-14   nfactor = {2.635202665e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.093364291e-06 wnfactor = -5.413638538e-06 pnfactor = 6.509329198e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.174890273e-04 leta0 = -3.498163991e-11 weta0 = 4.866968214e-11 peta0 = -9.734934157e-17   etab = -5.413834626e-04 letab = 5.984996690e-11 wetab = 8.677556799e-11 petab = -6.116640045e-17   dsub = -2.459730165e-01 ldsub = 1.560615841e-06 wdsub = 4.342425890e-07 pdsub = -1.975760454e-12   voffl = 0.0   minv = 0.0   pclm = -8.369341093e-01 lpclm = 1.378994291e-06 wpclm = 3.246299689e-06 ppclm = -4.563128340e-12   pdiblc1 = 0.39   pdiblc2 = 9.640714874e-03 lpdiblc2 = 6.283913268e-10 wpdiblc2 = -2.010988176e-08 ppdiblc2 = 2.873528573e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.422433131e-04 lalpha0 = -6.410195982e-11 walpha0 = 2.753629277e-10 palpha0 = -3.654057072e-16   alpha1 = 0.0   beta0 = 2.033543389e+01 lbeta0 = 1.519331398e-06 wbeta0 = 5.217087444e-06 pbeta0 = -8.254348308e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.985241777e-01 lkt1 = 3.523852532e-08 wkt1 = 1.654461724e-07 pkt1 = -1.710074717e-13   kt2 = 5.558860430e-02 lkt2 = -1.127332067e-07 wkt2 = -3.120821263e-07 pkt2 = 4.175396538e-13   at = 9.303874781e+04 lat = -2.423342765e-02 wat = -2.467999564e-01 pat = 2.710992505e-7   ute = -1.264284280e+00 lute = -5.859554146e-09 wute = -1.457558961e-07 pute = 6.231506525e-13   ua1 = 5.022996667e-09 lua1 = -3.613196855e-15 wua1 = -9.512251136e-15 pua1 = 1.326995007e-20   ub1 = -6.010179291e-18 lub1 = 5.169697097e-24 wub1 = 1.185747776e-23 pub1 = -1.832263935e-29   uc1 = -9.738967959e-11 luc1 = 1.567457371e-16 wuc1 = 2.279353881e-16 puc1 = -6.567060229e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.28 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.435192037e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.040314451e-08 wvth0 = -6.265890656e-09 pvth0 = 1.723248326e-14   k1 = 4.017951530e-01 lk1 = 3.068324389e-08 wk1 = 1.244930331e-07 pk1 = -1.092285213e-13   k2 = -1.278055775e-02 lk2 = -1.282594527e-08 wk2 = -1.856697009e-08 pk2 = 2.437596392e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -7.705737512e+04 lvsat = 1.449970086e-01 wvsat = 1.564806664e-01 pvsat = -1.266864132e-7   ua = -1.042312915e-09 lua = -5.535924573e-16 wua = -1.960187234e-15 pua = 2.277677291e-21   ub = 2.600433663e-18 lub = 2.840152221e-25 wub = 8.745150714e-25 pub = -1.971420410e-30   uc = 9.333316875e-11 luc = -1.328628834e-17 wuc = 1.562555000e-17 puc = -3.464438568e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.763993115e-02 lu0 = -6.120510191e-09 wu0 = -3.314281623e-08 pu0 = 2.074049259e-14   a0 = 2.915242744e+00 la0 = -8.520279092e-07 wa0 = -4.987705322e-06 pa0 = 3.361128926e-12   keta = -3.081660890e-01 lketa = 1.630079744e-07 wketa = -1.476930706e-07 pketa = 3.042797805e-14   a1 = 0.0   a2 = 0.38689047   ags = 4.855111323e+00 lags = -2.956199098e-06 wags = -4.757669466e-06 pags = 5.094379454e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.101075261e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.645020184e-09 wvoff = -3.191616171e-08 pvoff = 2.799366856e-14   nfactor = {1.447252242e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.482966187e-08 wnfactor = -3.693642387e-07 pnfactor = 1.464020823e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 9.798710349e-04 leta0 = -4.974583377e-10 weta0 = -1.691382690e-10 peta0 = 1.205032602e-16   etab = -9.533300678e-04 letab = 4.718810211e-10 wetab = 3.118884748e-10 petab = -2.863254554e-16   dsub = 1.628774799e+00 ldsub = -3.145162985e-07 wdsub = -3.082857690e-06 pdsub = 1.542060831e-12   voffl = 0.0   minv = 0.0   pclm = 5.663920943e-01 lpclm = -2.461959451e-08 wpclm = -1.982402633e-06 ppclm = 6.666458666e-13   pdiblc1 = 0.39   pdiblc2 = 1.215403446e-02 lpdiblc2 = -1.885443488e-09 wpdiblc2 = 9.865943438e-09 ppdiblc2 = -1.246684503e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.201471164e-05 lalpha0 = 5.615128849e-11 walpha0 = -1.082091522e-10 palpha0 = 1.824500508e-17   alpha1 = 0.0   beta0 = 1.948382264e+01 lbeta0 = 2.371117230e-06 wbeta0 = -4.677911575e-06 pbeta0 = 1.642679186e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.505104341e-01 lkt1 = -1.278506106e-08 wkt1 = -6.260637913e-08 pkt1 = 5.709183066e-14   kt2 = -6.591111411e-02 lkt2 = 8.791419133e-09 wkt2 = 1.425566021e-07 pkt2 = -3.719227559e-14   at = 1.189883417e+05 lat = -5.018834116e-02 wat = -1.065595145e-01 pat = 1.308300592e-7   ute = -2.224609197e+00 lute = 9.546622295e-07 wute = 4.528161239e-06 pute = -4.051724636e-12   ua1 = -2.672774255e-09 lua1 = 4.084151701e-15 wua1 = 2.265697420e-14 pua1 = -1.890586995e-20   ub1 = 4.515290151e-18 lub1 = -5.357930066e-24 wub1 = -3.078974708e-23 pub1 = 2.433332818e-29   uc1 = 1.828952524e-10 luc1 = -1.235966534e-16 wuc1 = -1.044527042e-15 puc1 = 6.160172621e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.29 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.987010887e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.800539931e-08 wvth0 = 4.536766225e-09 pvth0 = 1.182894028e-14   k1 = 3.087906387e-01 lk1 = 7.720456696e-08 wk1 = -1.086965420e-07 pk1 = 7.414070146e-15   k2 = 1.549311421e-02 lk2 = -2.696857736e-08 wk2 = 2.365218085e-08 pk2 = 3.257733526e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.647311091e+05 lvsat = -2.596730014e-02 wvsat = -2.304980492e-01 pvsat = 6.688227526e-8   ua = -3.279311410e-09 lua = 5.653653751e-16 wua = 8.777988285e-15 pua = -3.093611794e-21   ub = 4.580532150e-18 lub = -7.064399412e-25 wub = -8.610928914e-24 pub = 2.773246099e-30   uc = 5.023436147e-11 luc = 8.271950556e-18 wuc = -2.972766214e-18 puc = -2.534141492e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.330707724e-02 lu0 = 1.048855001e-09 wu0 = 5.221622986e-08 pu0 = -2.195652905e-14   a0 = 1.047946582e+00 la0 = 8.200296760e-08 wa0 = 3.118531796e-06 pa0 = -6.936514120e-13   keta = 7.400834395e-02 lketa = -2.815758786e-08 wketa = -1.892324881e-07 pketa = 5.120620239e-14   a1 = 0.0   a2 = 0.38689047   ags = -2.110592557e+00 lags = 5.280808107e-07 wags = 1.085827759e-05 pags = -2.716795345e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.252664425e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.937545596e-09 wvoff = 3.989233857e-08 pvoff = -7.925302320e-15   nfactor = {1.873418407e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.250431440e-07 wnfactor = 6.666204417e-06 pnfactor = -2.055205797e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.152977395e-03 leta0 = -1.584456896e-09 weta0 = -3.305146059e-08 peta0 = 1.656840530e-14   etab = 1.114097891e-01 letab = -5.573271298e-08 wetab = -2.708589624e-07 petab = 1.353546900e-13   dsub = 1.550686472e+00 ldsub = -2.754561269e-07 wdsub = 5.410655006e-07 pdsub = -2.706436687e-13   voffl = 0.0   minv = 0.0   pclm = 5.977801423e-01 lpclm = -4.032005308e-08 wpclm = -1.083194020e-06 ppclm = 2.168572223e-13   pdiblc1 = 0.39   pdiblc2 = 5.043193649e-03 lpdiblc2 = 1.671434639e-09 wpdiblc2 = -9.125198758e-10 ppdiblc2 = 4.144756738e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.333534370e-03 lalpha0 = 7.342037171e-10 walpha0 = -1.335533239e-09 palpha0 = 6.321586498e-16   alpha1 = 0.0   beta0 = 1.790638536e+01 lbeta0 = 3.160159243e-06 wbeta0 = -2.594495821e-06 pbeta0 = 6.005442088e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.436428223e-01 lkt1 = 3.380022519e-08 wkt1 = 2.851880441e-07 pkt1 = -1.168766788e-13   kt2 = -5.995567726e-02 lkt2 = 5.812479843e-09 wkt2 = 8.354506741e-08 pkt2 = -7.674410882e-15   at = -4.963579141e+01 lat = 9.355050347e-03 wat = 2.545761642e-01 pat = -4.981181295e-8   ute = -1.040825627e+00 lute = 3.625277688e-07 wute = -1.025221705e-06 pute = -1.273894720e-12   ua1 = 4.752237893e-09 lua1 = 3.701234990e-16 wua1 = -1.216202088e-14 pua1 = -1.489234522e-21   ub1 = -6.468664437e-18 lub1 = 1.362989385e-25 wub1 = 1.827583821e-23 pub1 = -2.095229143e-31   uc1 = -1.726173288e-10 luc1 = 5.423251729e-17 wuc1 = 5.907280504e-16 puc1 = -2.019455114e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.30 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.241865205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.940248175e-08 wvth0 = -2.137316466e-07 pvth0 = 6.644078851e-14   k1 = 3.530004470e-01 lk1 = 6.614305188e-08 wk1 = -7.530394912e-08 pk1 = -9.409235663e-16   k2 = 2.107949938e-03 lk2 = -2.361954233e-08 wk2 = 5.113554630e-08 pk2 = -3.618741925e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 9.824303140e+04 lvsat = 1.568884933e-02 wvsat = 1.968286641e-01 pvsat = -4.003700503e-8   ua = 3.273679703e-09 lua = -1.074225766e-15 wua = -1.608037877e-14 pua = 3.126075936e-21   ub = -1.755483646e-18 lub = 8.788628910e-25 wub = 1.263461164e-23 pub = -2.542494374e-30   uc = 2.180341589e-10 luc = -3.371239775e-17 wuc = -4.329143169e-16 puc = 8.223211077e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 6.268115081e-02 lu0 = -8.802735076e-09 wu0 = -1.467920090e-07 pu0 = 2.783632735e-14   a0 = 4.917206317e+00 la0 = -8.861051644e-07 wa0 = 1.237440515e-06 pa0 = -2.229929680e-13   keta = -2.059196544e-02 lketa = -4.488117449e-09 wketa = 5.461917087e-07 pketa = -1.328006088e-13   a1 = 0.0   a2 = 0.38689047   ags = -3.258300685e+00 lags = 8.152431229e-07 wags = 9.311917680e-07 pags = -2.329888363e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.811757498e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.692633382e-08 wvoff = 6.812998134e-08 pvoff = -1.499050173e-14   nfactor = {3.231126385e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.652696782e-08 wnfactor = -6.701689696e-06 pnfactor = 1.289508150e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.080279028e-05 lcit = -1.451887142e-12 wcit = -1.690329598e-11 pcit = 4.229289171e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.862125449e-01 leta0 = 7.081624352e-08 weta0 = 3.179233417e-07 peta0 = -7.124724511e-14   etab = -3.460130104e-01 letab = 5.871675856e-08 wetab = 9.252439352e-07 petab = -1.639162355e-13   dsub = 8.547825480e-01 ldsub = -1.013374855e-07 wdsub = -2.254823739e-06 pdsub = 4.289017985e-13   voffl = 0.0   minv = 0.0   pclm = 1.486509040e+00 lpclm = -2.626844669e-07 wpclm = -2.142096535e-06 ppclm = 4.817999260e-13   pdiblc1 = -1.191545093e+00 lpdiblc1 = 3.957104899e-07 wpdiblc1 = 5.486899685e-08 ppdiblc1 = -1.372849736e-14   pdiblc2 = 2.401123381e-02 lpdiblc2 = -3.074463850e-09 wpdiblc2 = 1.572682752e-08 ppdiblc2 = -1.849117749e-17   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.581651483e-03 lalpha0 = 7.962838593e-10 walpha0 = 2.144749002e-08 palpha0 = -5.068267686e-15   alpha1 = 0.0   beta0 = 2.435523583e+01 lbeta0 = 1.546624611e-06 wbeta0 = 3.146638076e-05 pbeta0 = -7.921657417e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 7.438810179e-02 lkt1 = -7.079320218e-08 wkt1 = -7.702123340e-07 pkt1 = 1.471897728e-13   kt2 = -1.565831085e-02 lkt2 = -5.270942718e-09 wkt2 = 1.597594913e-08 pkt2 = 9.231720359e-15   at = -1.277681424e+05 lat = 4.131085928e-02 wat = 4.310543651e-01 pat = -9.396754118e-8   ute = 5.041109255e+00 lute = -1.159202748e-06 wute = -1.937243607e-05 pute = 3.316670050e-12   ua1 = 2.035236894e-08 lua1 = -3.533107289e-15 wua1 = -5.896274517e-14 pua1 = 1.022054070e-20   ub1 = -1.922887503e-17 lub1 = 3.328967431e-24 wub1 = 5.493357185e-23 pub1 = -9.381471160e-30   uc1 = 1.352286275e-10 luc1 = -2.279208018e-17 wuc1 = -6.630205513e-16 puc1 = 1.117486575e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.31 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.227389161e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.365903353e-08 wvth0 = 8.989836799e-07 pvth0 = -1.340760769e-13   k1 = 6.373641371e-01 lk1 = 1.489929310e-08 wk1 = 8.045236970e-07 pk1 = -1.594902645e-13   k2 = -6.338624952e-02 lk2 = -1.181716012e-08 wk2 = -3.660894222e-07 pk2 = 7.156728352e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.239534837e+05 lvsat = -6.964802732e-03 wvsat = -1.744209976e-01 pvsat = 2.686404025e-8   ua = -2.811561021e-09 lua = 2.236503841e-17 wua = 3.510164699e-15 pua = -4.042379505e-22   ub = 1.192927979e-18 lub = 3.475443741e-25 wub = 3.729821348e-24 pub = -9.378066407e-31   uc = 1.351327949e-10 luc = -1.877315746e-17 wuc = -1.168309304e-16 puc = 2.527230410e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.673595471e-02 lu0 = 5.508624424e-09 wu0 = 1.304087248e-07 pu0 = -2.211663089e-14   a0 = 0.0   keta = -3.157490865e-01 lketa = 4.870067156e-08 wketa = 1.543545613e-06 pketa = -3.125287690e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.302900042e+00 lags = -6.708054177e-09 wags = -2.014672151e-06 pags = 2.978705712e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {2.446887271e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.981657423e-08 wvoff = -1.128596822e-06 pvoff = 2.006656518e-13   nfactor = {4.677840638e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.972321098e-07 wnfactor = -1.179181111e-05 pnfactor = 2.206773479e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.810514402e-05 lcit = -4.569857797e-12 wcit = -1.402278864e-10 pcit = 2.645299700e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.648820147e-01 leta0 = -6.453475158e-08 weta0 = -1.105489358e-06 peta0 = 1.852588404e-13   etab = 2.487336950e-02 letab = -8.118821532e-09 wetab = -3.316443884e-07 petab = 6.258132487e-14   dsub = 4.548434513e-01 ldsub = -2.926646061e-08 wdsub = 7.523762199e-07 pdsub = -1.130106701e-13   voffl = 0.0   minv = 0.0   pclm = -1.907269132e+00 lpclm = 3.488913285e-07 wpclm = 6.802329074e-06 ppclm = -1.130030291e-12   pdiblc1 = 2.415904892e+00 lpdiblc1 = -2.543700346e-07 wpdiblc1 = -4.176463378e-06 ppdiblc1 = 7.487787533e-13   pdiblc2 = 4.836053998e-02 lpdiblc2 = -7.462330567e-09 wpdiblc2 = -1.048886381e-08 ppdiblc2 = 4.705707480e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.151622438e-02 lalpha0 = -1.564018860e-09 walpha0 = -2.889034167e-08 palpha0 = 4.002861275e-15   alpha1 = 0.0   beta0 = 4.296945561e+01 lbeta0 = -1.807750864e-06 wbeta0 = -3.171248488e-05 pbeta0 = 3.463490066e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.111787218e+00 lkt1 = 1.429615213e-07 wkt1 = 3.134727624e-06 pkt1 = -5.564999323e-13   kt2 = -2.077739399e-01 lkt2 = 2.934925421e-08 wkt2 = 3.930524762e-07 pkt2 = -5.871935521e-14   at = 3.290714399e+05 lat = -4.101391764e-02 wat = -9.961046364e-01 pat = 1.632136467e-7   ute = -2.982586278e+00 lute = 2.867073052e-07 wute = 2.787627648e-06 pute = -6.766842324e-13   ua1 = -8.385726141e-10 lua1 = 2.856063334e-16 wua1 = -2.243474255e-16 pua1 = -3.644122666e-22   ub1 = 6.081348890e-19 lub1 = -2.457609423e-25 wub1 = 3.426778753e-24 pub1 = -9.968950964e-32   uc1 = 8.366629439e-11 luc1 = -1.350028995e-17 wuc1 = 2.235265100e-16 puc1 = -4.801155572e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.32 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.426083+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.50407   k2 = -0.048504361   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169790.0   ua = -1.10059665e-9   ub = 2.406442e-18   uc = 6.9010287e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03195911   a0 = 1.687182   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.523358   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.40896304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0067115   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.8823913e-5   alpha1 = 0.0   beta0 = 17.79575   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.2558   kt2 = -0.03478   at = 318480.0   ute = -1.261   ua1 = 2.0849e-9   ub1 = -2.0887e-18   uc1 = -4.6822e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.33 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.426083+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.50407   k2 = -0.048504361   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169790.0   ua = -1.10059665e-9   ub = 2.406442e-18   uc = 6.9010287e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03195911   a0 = 1.687182   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.523358   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.40896304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0067115   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.8823913e-5   alpha1 = 0.0   beta0 = 17.79575   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.2558   kt2 = -0.03478   at = 318480.0   ute = -1.261   ua1 = 2.0849e-9   ub1 = -2.0887e-18   uc1 = -4.6822e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.34 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.171711866e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.564908039e-8   k1 = 5.656663130e-01 lk1 = -2.463978791e-7   k2 = -7.777382181e-02 lk2 = 1.170838435e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.014804969e+05 lvsat = -5.267889841e-1   ua = -9.669357012e-10 lua = -5.346711959e-16   ub = 2.266329640e-18 lub = 5.604781632e-25   uc = 4.910553397e-11 luc = 7.962309259e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.220115181e-02 lu0 = -9.682168455e-10   a0 = 1.569670956e+00 la0 = 4.700682644e-7   keta = 2.518358105e-01 lketa = -1.007394868e-6   a1 = 0.0   a2 = 0.38689047   ags = -6.708863975e-01 lags = 4.777222410e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.117054424e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.239610567e-8   nfactor = {1.470631910e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.466881238e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081487e-01 leta0 = -3.180488942e-7   etab = -1.395149546e-01 letab = 2.780740688e-7   dsub = 7.757925865e-01 ldsub = -8.632145834e-7   voffl = 0.0   minv = 0.0   pclm = 2.162416646e-01 lpclm = -6.496998794e-8   pdiblc1 = 0.39   pdiblc2 = 5.439769661e-03 lpdiblc2 = 5.087182061e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.437439074e-05 lalpha0 = 4.128143706e-10   alpha1 = 0.0   beta0 = 1.412179646e+01 lbeta0 = 1.469656733e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.581402399e-01 lkt1 = 9.361439149e-9   kt2 = -3.331384973e-02 lkt2 = -5.864901621e-9   at = 5.942612647e+05 lat = -1.103181594e+0   ute = -1.311705197e+00 lute = 2.028311816e-7   ua1 = 1.941185271e-09 lua1 = 5.748883785e-16   ub1 = -1.677657873e-18 lub1 = -1.644252774e-24   uc1 = -4.015731694e-11 luc1 = -2.666009850e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.35 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.331056750e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.776837100e-9   k1 = 4.472409758e-01 lk1 = -9.522927600e-9   k2 = -1.486350343e-02 lk2 = -8.749689886e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.929206970e+03 lvsat = 8.009262259e-2   ua = -9.814760732e-10 lua = -5.055874710e-16   ub = 2.585118907e-18 lub = -7.716572279e-26   uc = 1.043061550e-10 luc = -3.078946550e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.617351938e-02 lu0 = -8.913766328e-9   a0 = 2.104663484e+00 la0 = -6.000264640e-7   keta = -3.181836038e-01 lketa = 1.327608142e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.420149060e+00 lags = 5.947228335e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.197059596e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.606568755e-9   nfactor = {7.767361783e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.141245589e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.341970090e-04 leta0 = -6.840102829e-11   etab = -5.115939811e-04 letab = 3.885194412e-11   dsub = -9.690039310e-02 ldsub = 8.823502778e-7   voffl = 0.0   minv = 0.0   pclm = 2.774992126e-01 lpclm = -1.874976417e-7   pdiblc1 = 0.39   pdiblc2 = 2.737124795e-03 lpdiblc2 = 1.049302583e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.367735942e-04 lalpha0 = -1.895433346e-10   alpha1 = 0.0   beta0 = 2.212642568e+01 lbeta0 = -1.314332060e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.417275954e-01 lkt1 = -2.346721444e-8   kt2 = -5.154713609e-02 lkt2 = 3.060540891e-8   at = 8.313946770e+03 lat = 6.883316114e-2   ute = -1.314321320e+00 lute = 2.080639644e-7   ua1 = 1.757503445e-09 lua1 = 9.422896848e-16   ub1 = -1.939585200e-18 lub1 = -1.120344424e-24   uc1 = -1.914096071e-11 luc1 = -6.869711931e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.36 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.413681647e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.487346399e-9   k1 = 4.445327921e-01 lk1 = -6.814188722e-9   k2 = -1.915447641e-02 lk2 = -4.457837259e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.333859204e+04 lvsat = 1.015063966e-1   ua = -1.715232293e-09 lua = 2.283191692e-16   ub = 2.900648933e-18 lub = -3.927604322e-25   uc = 9.869731724e-11 luc = -2.517947798e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.626222043e-02 lu0 = 9.995644382e-10   a0 = 1.202996328e+00 la0 = 3.018255340e-7   keta = -3.588681483e-01 lketa = 1.734536990e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.221834702e+00 lags = -1.207332154e-06 pags = 2.067951531e-25   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.210641344e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.965022029e-9   nfactor = {1.320451929e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.974183766e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 9.218068821e-04 leta0 = -4.560903615e-10   etab = -8.462608067e-04 letab = 3.735873764e-10   dsub = 5.704500403e-01 ldsub = 2.148630376e-7   voffl = 0.0   minv = 0.0   pclm = -1.141536851e-01 lpclm = 2.042355448e-7   pdiblc1 = 0.39   pdiblc2 = 1.554094792e-02 lpdiblc2 = -2.313422074e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.513277829e-05 lalpha0 = 6.241467867e-11   alpha1 = 0.0   beta0 = 1.787792637e+01 lbeta0 = 2.935038185e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.720027921e-01 lkt1 = 6.814188722e-9   kt2 = -1.697237066e-02 lkt2 = -3.976444344e-9   at = 8.240716152e+04 lat = -5.275242723e-3   ute = -6.701212400e-01 lute = -4.362681766e-7   ua1 = 5.105215898e-09 lua1 = -2.406109050e-15   ub1 = -6.054627417e-18 lub1 = 2.995541377e-24   uc1 = -1.756840078e-10 luc1 = 8.787801914e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.37 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.002585307e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.394460195e-8   k1 = 2.714758311e-01 lk1 = 7.974976846e-8   k2 = 2.361275226e-02 lk2 = -2.585021888e-08 pk2 = 1.615587134e-27   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.856026455e+05 lvsat = -3.007055143e-3   ua = -2.658857929e-10 lua = -4.966511971e-16   ub = 1.624456916e-18 lub = 2.455971958e-25   uc = 4.921383039e-11 luc = -4.275904335e-19   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.123256535e-02 lu0 = -6.488676944e-9   a0 = 2.118518027e+00 la0 = -1.561229977e-7   keta = 9.046075971e-03 lketa = -1.057883553e-8   a1 = 0.0   a2 = 0.38689047   ags = 1.616982691e+00 lags = -4.045771543e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.115716652e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.168414601e-10   nfactor = {2.475805952e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.950451763e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -8.193371853e-03 leta0 = 4.103367618e-09 weta0 = 3.374896899e-22 peta0 = -1.901154782e-28   etab = 1.842568958e-02 letab = -9.266338567e-09 wetab = 1.588186776e-22 petab = 1.956375045e-28   dsub = 1.736430698e+00 ldsub = -3.683663175e-7   voffl = 0.0   minv = 0.0   pclm = 2.259267628e-01 lpclm = 3.412560437e-8   pdiblc1 = 0.39   pdiblc2 = 4.729931580e-03 lpdiblc2 = 3.094302354e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.792014143e-03 lalpha0 = 9.512196218e-10 walpha0 = -7.940933881e-23 palpha0 = -3.786532345e-29   alpha1 = 0.0   beta0 = 1.701571202e+01 lbeta0 = 3.366322119e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.457396434e-01 lkt1 = -6.322769573e-9   kt2 = -3.127520536e-02 lkt2 = 3.177905087e-9   at = 8.734468622e+04 lat = -7.745017266e-03 wat = -1.421085472e-14   ute = -1.392777492e+00 lute = -7.479190611e-8   ua1 = 5.770961539e-10 lua1 = -1.411209128e-16   ub1 = -1.946894389e-19 lub1 = 6.437110077e-26 pub1 = 5.605193857e-45   uc1 = 3.017572382e-11 luc1 = -1.509404793e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.38 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.508138526e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.659379626e-8   k1 = 3.271490968e-01 lk1 = 6.582003901e-8   k2 = 1.966244650e-02 lk2 = -2.486183262e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.658130166e+05 lvsat = 1.944408958e-3   ua = -2.246608517e-09 lua = -1.064467802e-18   ub = 2.581895389e-18 lub = 6.041302438e-27   uc = 6.941752254e-11 luc = -5.482655230e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.228842004e-02 lu0 = 7.532929330e-10   a0 = 5.342011503e+00 la0 = -9.626571829e-7   keta = 1.669120541e-01 lketa = -5.007769258e-08 pketa = 3.231174268e-27   a1 = 0.0   a2 = 0.38689047   ags = -2.938628679e+00 lags = 7.352595885e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.577871755e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.178019322e-8   nfactor = {9.304804108e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.061526946e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.770715537e-01 leta0 = 4.635753310e-08 weta0 = -6.776263578e-21 peta0 = -1.615587134e-27   etab = -2.838285576e-02 letab = 2.445393521e-9   dsub = 8.071639565e-02 ldsub = 4.590167963e-8   voffl = 0.0   minv = 0.0   pclm = 7.511413951e-01 lpclm = -9.728572270e-8   pdiblc1 = -1.172708927e+00 lpdiblc1 = 3.909975871e-7   pdiblc2 = 2.941015021e-02 lpdiblc2 = -3.080811749e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 5.781130712e-03 lalpha0 = -9.436190868e-10   alpha1 = 0.0   beta0 = 3.515743729e+01 lbeta0 = -1.172828254e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.900207243e-01 lkt1 = -2.026392173e-8   kt2 = -1.017387264e-02 lkt2 = -2.101753865e-9   at = 2.020998471e+04 lat = 9.052420725e-3   ute = -1.609320571e+00 lute = -2.061174493e-8   ua1 = 1.108465099e-10 lua1 = -2.446292064e-17 wua1 = -6.310887242e-30 pua1 = -1.504632769e-36   ub1 = -3.705412919e-19 lub1 = 1.083701136e-25 pub1 = -5.605193857e-45   uc1 = -9.238196496e-11 luc1 = 1.557049859e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.39 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-2.747837204e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.478396174e-07 wvth0 = 9.055595297e-06 pvth0 = -1.631863550e-12   k1 = 9.135518283e-01 lk1 = -3.985266522e-8   k2 = 9.053958189e-01 lk2 = -1.844754150e-07 wk2 = -3.188112836e-06 pk2 = 5.745138736e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.319511609e+06 lvsat = -9.267778459e-01 wvsat = -1.501757799e+01 pvsat = 2.706242642e-6   ua = 3.400725040e-09 lua = -1.018742211e-15 wua = -1.458597611e-14 pua = 2.628465824e-21   ub = 1.280747794e-17 lub = -1.836659800e-24 wub = -3.010289809e-23 pub = 5.424692751e-30   uc = 9.502550528e-11 luc = -1.009734176e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -9.030821675e-03 lu0 = 4.595126887e-09 wu0 = 1.079639805e-07 pu0 = -1.945564911e-14   a0 = 0.0   keta = 2.141399654e-01 lketa = -5.858839834e-8   a1 = 0.0   a2 = 0.38689047   ags = 6.112763500e-01 lags = 9.554895285e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.427511353e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.070623598e-9   nfactor = {-7.465962963e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.402786847e-05 wnfactor = 2.193150663e-04 pnfactor = -3.952167152e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.003416667e-05 lcit = 4.511282004e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.537479252e-02 leta0 = -9.366107155e-10   etab = -8.897796674e-02 letab = 1.336493549e-8   dsub = 7.131292568e-01 ldsub = -6.806228002e-8   voffl = 0.0   minv = 0.0   pclm = 4.279256783e-01 lpclm = -3.904063446e-8   pdiblc1 = 9.821524968e-01 lpdiblc1 = 2.680784218e-9   pdiblc2 = 4.475978205e-02 lpdiblc2 = -5.846892154e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.598360187e-03 lalpha0 = -1.898629242e-10   alpha1 = 0.0   beta0 = 3.208276822e+01 lbeta0 = -6.187575149e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.565585167e-02 lkt1 = -4.808124360e-8   kt2 = -7.284161117e-02 lkt2 = 9.191285955e-9   at = -1.288472717e+04 lat = 1.501625328e-2   ute = -2.025612050e+00 lute = 5.440606097e-8   ua1 = -9.155896090e-10 lua1 = 1.605060002e-16 wua1 = -2.524354897e-29   ub1 = 1.784525486e-18 lub1 = -2.799836950e-25 wub1 = -1.880790961e-37   uc1 = 1.604014744e-10 luc1 = -2.998234110e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.40 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.315918668e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.599201989e-8   k1 = 4.704915538e-01 wk1 = 9.747688625e-8   k2 = -3.826178801e-02 wk2 = -2.973377968e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.344055188e+05 wvsat = 1.027197335e-1   ua = -1.242306378e-09 wua = 4.113776724e-16   ub = 2.698049927e-18 wub = -8.465261471e-25   uc = 1.226848409e-10 wuc = -1.558150829e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.580758645e-02 wu0 = -1.117197320e-8   a0 = 1.420322159e+00 wa0 = 7.746834445e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.837023036e-01 wags = 1.151189003e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.200616203e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.526176139e-8   nfactor = {9.082464495e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.453560234e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -7.517037037e-07 wcit = 1.669696578e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 5.724967781e-03 wpdiblc2 = 2.863863571e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.547524350e-05 walpha0 = 9.721053625e-12   alpha1 = 0.0   beta0 = 1.779849586e+01 wbeta0 = -7.971131465e-9   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.536948764e-01 wkt1 = -6.111089477e-9   kt2 = -3.295786027e-02 wkt2 = -5.289598760e-9   at = 6.178561778e+05 wat = -8.690770690e-1   ute = -1.353257327e+00 wute = 2.678193312e-7   ua1 = 2.224436332e-09 wua1 = -4.050683899e-16   ub1 = -2.805017179e-18 wub1 = 2.079440119e-24   uc1 = -1.736355633e-10 wuc1 = 3.681347016e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.41 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.315918668e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.599201989e-8   k1 = 4.704915538e-01 wk1 = 9.747688625e-8   k2 = -3.826178801e-02 wk2 = -2.973377968e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.344055188e+05 wvsat = 1.027197335e-1   ua = -1.242306378e-09 wua = 4.113776724e-16   ub = 2.698049927e-18 wub = -8.465261471e-25   uc = 1.226848409e-10 wuc = -1.558150829e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.580758645e-02 wu0 = -1.117197320e-8   a0 = 1.420322159e+00 wa0 = 7.746834445e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.837023036e-01 wags = 1.151189003e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.200616203e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.526176139e-8   nfactor = {9.082464495e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.453560234e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -7.517037037e-07 wcit = 1.669696578e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 5.724967781e-03 wpdiblc2 = 2.863863571e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.547524350e-05 walpha0 = 9.721053625e-12   alpha1 = 0.0   beta0 = 1.779849586e+01 wbeta0 = -7.971131465e-9   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.536948764e-01 wkt1 = -6.111089477e-9   kt2 = -3.295786027e-02 wkt2 = -5.289598760e-9   at = 6.178561778e+05 wat = -8.690770690e-1   ute = -1.353257327e+00 wute = 2.678193312e-7   ua1 = 2.224436332e-09 wua1 = -4.050683899e-16   ub1 = -2.805017179e-18 wub1 = 2.079440119e-24   uc1 = -1.736355633e-10 wuc1 = 3.681347016e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.42 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.291106571e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.925347422e-09 wvth0 = -3.465980513e-08 pvth0 = 7.467496786e-14   k1 = 5.162805649e-01 lk1 = -1.831654312e-07 wk1 = 1.433648513e-07 pk1 = -1.835612671e-13   k2 = -6.748091971e-02 lk2 = 1.168825167e-07 wk2 = -2.987988309e-08 pk2 = 5.844435772e-16   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.359827605e+05 lvsat = -4.063297902e-01 wvsat = 1.901373088e-01 pvsat = -3.496882216e-7   ua = -1.102473391e-09 lua = -5.593606135e-16 wua = 3.934604927e-16 pua = 7.167239182e-23   ub = 2.570700525e-18 lub = 5.094237141e-25 wub = -8.835765041e-25 pub = 1.482090236e-31   uc = 1.133777678e-10 luc = 3.723020025e-17 wuc = -1.865797239e-16 puc = 1.230648707e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.644552064e-02 lu0 = -2.551867521e-09 wu0 = -1.232123294e-08 pu0 = 4.597274566e-15   a0 = 1.060620817e+00 la0 = 1.438879107e-06 wa0 = 1.477752193e-06 pa0 = -2.812419124e-12   keta = 3.330351821e-01 lketa = -1.332209001e-06 wketa = -2.357185277e-07 pketa = 9.429224330e-13   a1 = 0.0   a2 = 0.38689047   ags = -1.121098219e+00 lags = 6.419531076e-06 wags = 1.306946910e-06 pags = -4.767556365e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.212276524e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.664367742e-09 wvoff = 2.764259485e-08 pvoff = -4.952587190e-14   nfactor = {4.878903101e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.681510731e-06 wnfactor = 2.852859556e-06 pnfactor = -5.597484146e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -7.517037037e-07 wcit = 1.669696578e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081487e-01 leta0 = -3.180488942e-7   etab = -1.395239626e-01 letab = 2.781101030e-07 wetab = 2.615012853e-11 petab = -1.046058749e-16   dsub = 8.425347769e-01 ldsub = -1.130197027e-06 wdsub = -1.937499092e-07 pdsub = 7.750393555e-13   voffl = 0.0   minv = 0.0   pclm = 2.746504503e-01 lpclm = -2.986171045e-07 wpclm = -1.695583685e-07 ppclm = 6.782682335e-13   pdiblc1 = 0.39   pdiblc2 = 7.797965877e-03 lpdiblc2 = -8.292417349e-09 wpdiblc2 = -6.845749287e-09 ppdiblc2 = 3.884044190e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -9.129340858e-05 lalpha0 = 5.071005959e-10 walpha0 = 7.814483203e-11 palpha0 = -2.737091405e-16   alpha1 = 0.0   beta0 = 1.380735512e+01 lbeta0 = 1.596538116e-05 wbeta0 = 9.128106293e-07 pbeta0 = -3.683315803e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.712556842e-01 lkt1 = 7.024683116e-08 wkt1 = 3.807361045e-08 pkt1 = -1.767478576e-13   kt2 = -3.063922014e-02 lkt2 = -9.275035822e-09 wkt2 = -7.764342725e-09 pkt2 = 9.899483180e-15   at = 1.200459012e+06 lat = -2.330530772e+00 wat = -1.759767813e+00 pat = 3.562945569e-6   ute = -1.391997754e+00 lute = 1.549696489e-07 wute = 2.330860825e-07 pute = 1.389401148e-13   ua1 = 2.010543625e-09 lua1 = 8.556146758e-16 wua1 = -2.013445278e-16 pua1 = -8.149372119e-22   ub1 = -2.413877986e-18 lub1 = -1.564636955e-24 wub1 = 2.137217542e-24 pub1 = -2.311215371e-31   uc1 = -2.428368405e-10 luc1 = 2.768192952e-16 wuc1 = 5.883705497e-16 puc1 = -8.809885409e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.43 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.353166530e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.487916554e-09 wvth0 = -6.418380579e-09 pvth0 = 1.818632927e-14   k1 = 4.344271963e-01 lk1 = -1.944191414e-08 wk1 = 3.719788925e-08 pk1 = 2.879442118e-14   k2 = -4.404205582e-03 lk2 = -9.283842271e-09 wk2 = -3.036292329e-08 pk2 = 1.550623006e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -5.634132838e+03 lvsat = 7.695352801e-02 wvsat = 1.075525160e-02 pvsat = 9.112666006e-9   ua = -1.301740131e-09 lua = -1.607862843e-16 wua = 9.297137490e-16 pua = -1.000944053e-21   ub = 2.979579834e-18 lub = -3.084187241e-25 wub = -1.145104292e-24 pub = 6.713182128e-31   uc = 1.571156916e-10 luc = -5.025461357e-17 wuc = -1.533039724e-16 puc = 5.650654625e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.911956012e-02 lu0 = -7.900494674e-09 wu0 = -8.552238440e-09 pu0 = -2.941487081e-15   a0 = 1.994022201e+00 la0 = -4.281150079e-07 wa0 = 3.211872194e-07 pa0 = -4.990520807e-13   keta = -3.966592926e-01 lketa = 1.273295362e-07 wketa = 2.278117856e-07 pketa = 1.576678283e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.762001376e+00 lags = 6.527408500e-07 wags = -9.923836002e-07 pags = -1.684239810e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.205988796e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.406693121e-09 wvoff = 2.592111089e-09 pvoff = 5.802309697e-16   nfactor = {9.468728768e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.634515058e-07 wnfactor = -4.939000302e-07 pnfactor = 1.096721112e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.504586507e-06 lcit = 1.150694495e-11 wcit = 3.339735445e-11 pcit = -3.340420090e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.969988687e-04 leta0 = 6.002877740e-12 weta0 = 1.079847131e-10 peta0 = -2.159915630e-16   etab = -4.926113143e-04 letab = 1.889890158e-11 wetab = -5.510592236e-11 petab = 5.792288437e-17   dsub = -4.749252902e-01 ldsub = 1.504993186e-06 wdsub = 1.097391155e-06 pdsub = -1.807507457e-12   voffl = 0.0   minv = 0.0   pclm = 3.009139124e-01 lpclm = -3.511494128e-07 wpclm = -6.797193698e-08 ppclm = 4.750745452e-13   pdiblc1 = 0.39   pdiblc2 = -4.240004091e-03 lpdiblc2 = 1.578599037e-08 wpdiblc2 = 2.025432607e-08 ppdiblc2 = -1.536526433e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.769740897e-04 lalpha0 = -2.295098956e-10 walpha0 = -1.167004305e-10 palpha0 = 1.160213279e-16   alpha1 = 0.0   beta0 = 2.272093434e+01 lbeta0 = -1.863604571e-06 wbeta0 = -1.725834874e-06 pbeta0 = 1.594516126e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.120692831e-01 lkt1 = -4.813810441e-08 wkt1 = -8.609689423e-08 pkt1 = 7.161860674e-14   kt2 = -5.163938101e-02 lkt2 = 3.272959095e-08 wkt2 = 2.677833158e-10 pkt2 = -6.166415487e-15   at = -4.881646521e+03 lat = 8.039764081e-02 wat = 3.830627950e-02 pat = -3.357122191e-8   ute = -1.507366702e+00 lute = 3.857311944e-07 wute = 5.604030209e-07 pute = -5.157608619e-13   ua1 = 1.366954770e-09 lua1 = 2.142924321e-15 wua1 = 1.133747180e-15 pua1 = -3.485394322e-21   ub1 = -1.797576345e-18 lub1 = -2.797366580e-24 wub1 = -4.122460265e-25 pub1 = 4.868328240e-30   uc1 = -7.749328078e-11 luc1 = -5.390171964e-17 wuc1 = 1.693944511e-16 puc1 = -4.295045344e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.44 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.332302752e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.011111317e-10 wvth0 = 2.362396754e-08 pvth0 = -1.186217753e-14   k1 = 4.473731102e-01 lk1 = -3.239048188e-08 wk1 = -8.245329705e-09 pk1 = 7.424695599e-14   k2 = -1.318027684e-02 lk2 = -5.059719173e-10 wk2 = -1.734286238e-08 pk2 = -1.147210701e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3.063193675e+04 lvsat = 1.019564565e-01 wvsat = 2.117228795e-02 pvsat = -1.306505841e-9   ua = -2.348131754e-09 lua = 8.858198493e-16 wua = 1.837281819e-15 pua = -1.908698175e-21   ub = 3.582816030e-18 lub = -9.117785838e-25 wub = -1.980303797e-24 pub = 1.506688934e-30   uc = 1.750756877e-10 luc = -6.821829147e-17 wuc = -2.217233542e-16 puc = 1.249399540e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.526540918e-02 lu0 = 5.956496377e-09 wu0 = 2.893703201e-09 pu0 = -1.438977514e-14   a0 = 3.722964321e-01 la0 = 1.193943214e-06 wa0 = 2.411488569e-06 pa0 = -2.589781942e-12   keta = -5.127860622e-01 lketa = 2.434801117e-07 wketa = 4.468175473e-07 pketa = -2.032838751e-13   a1 = 0.0   a2 = 0.38689047   ags = 3.352322489e+00 lags = -9.379062794e-07 wags = -3.788008279e-07 pags = -7.821325377e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.367034453e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.951456026e-08 wvoff = 4.540029390e-08 pvoff = -4.223672752e-14   nfactor = {4.610889690e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.249334999e-06 wnfactor = 2.494696298e-06 pnfactor = -1.892487879e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.103579914e-03 leta0 = -3.601317517e-09 weta0 = -9.236559841e-09 peta0 = 9.130468623e-15   etab = -8.776634680e-04 letab = 4.040299910e-10 wetab = 9.116066977e-11 petab = -8.837369241e-17   dsub = 1.059531073e+00 ldsub = -2.977774020e-08 wdsub = -1.419782674e-06 pdsub = 7.101823923e-13   voffl = 0.0   minv = 0.0   pclm = -3.592882874e-01 lpclm = 3.091881285e-07 wpclm = 7.116159452e-07 ppclm = -3.046731524e-13   pdiblc1 = 0.39   pdiblc2 = 8.060898074e-03 lpdiblc2 = 3.482566520e-09 wpdiblc2 = 2.171428550e-08 ppdiblc2 = -1.682552305e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.124854138e-05 lalpha0 = 2.626807649e-11 walpha0 = -1.056135157e-10 palpha0 = 1.049321403e-16   alpha1 = 0.0   beta0 = 1.858874848e+01 lbeta0 = 2.269428393e-06 wbeta0 = -2.063488132e-06 pbeta0 = 1.932238603e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.761707798e-01 lkt1 = 1.597653317e-08 wkt1 = 1.209950167e-08 pkt1 = -2.659791943e-14   kt2 = -2.542361889e-02 lkt2 = 6.508454593e-09 wkt2 = 2.453363555e-08 pkt2 = -3.043724222e-14   at = 9.011252014e+04 lat = -1.461599965e-02 wat = -2.236834785e-02 pat = 2.711584374e-8   ute = -2.255560975e-01 lute = -8.963421809e-07 wute = -1.290554826e-06 pute = 1.335576432e-12   ua1 = 8.066994374e-09 lua1 = -4.558488792e-15 wua1 = -8.597924445e-15 pua1 = 6.248272296e-21   ub1 = -1.053560686e-17 lub1 = 5.942455227e-24 wub1 = 1.300810407e-23 pub1 = -8.554773030e-30   uc1 = -2.762931828e-10 luc1 = 1.449389364e-16 wuc1 = 2.920644106e-16 puc1 = -1.656455603e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.45 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.977348100e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.266660193e-08 wvth0 = 7.326260453e-09 pvth0 = -3.709982958e-15   k1 = 1.867077735e-01 lk1 = 9.799562284e-08 wk1 = 2.460782805e-07 pk1 = -5.296698545e-14   k2 = 5.508046195e-02 lk2 = -3.465033477e-08 wk2 = -9.134950252e-08 pk2 = 2.554638442e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.461036724e+05 lvsat = 1.355242108e-02 wvsat = 1.146639389e-01 pvsat = -4.807149708e-8   ua = 1.129877140e-09 lua = -8.538975895e-16 wua = -4.051843963e-15 pua = 1.037071987e-21   ub = 5.606386643e-19 lub = 5.999296455e-25 wub = 3.088221831e-24 pub = -1.028612928e-30   uc = 2.334215879e-11 luc = 7.679578339e-18 wuc = 7.510442777e-17 puc = -2.353478666e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 5.593410394e-02 lu0 = -9.384138089e-09 wu0 = -4.267797846e-08 pu0 = 8.405407884e-15   a0 = 4.048120318e+00 la0 = -6.447222723e-07 wa0 = -5.601558266e-06 pa0 = 1.418384150e-12   keta = -1.175502637e-02 lketa = -7.138117525e-09 wketa = 6.038476804e-08 pketa = -9.988266742e-15   a1 = 0.0   a2 = 0.38689047   ags = 2.955768766e+00 lags = -7.395481241e-07 wags = -3.886442423e-06 pags = 9.724073265e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.572350632e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.985860106e-09 wvoff = -7.503617126e-08 pvoff = 1.800619454e-14   nfactor = {3.405443284e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.234457511e-07 wnfactor = -2.698699991e-06 pnfactor = 7.052749121e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.075642010e-05 lcit = -2.879390116e-12 wcit = -1.671065730e-11 pcit = 8.358754333e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.055327524e-02 leta0 = 8.732164716e-09 weta0 = 3.588030514e-08 peta0 = -1.343721282e-14   etab = 3.000010687e-02 letab = -1.504118512e-08 wetab = -3.360007043e-08 petab = 1.676414856e-14   dsub = 1.834504877e+00 ldsub = -4.174235120e-07 wdsub = -2.847054173e-07 pdsub = 1.424110733e-13   voffl = 0.0   minv = 0.0   pclm = 3.814512036e-01 lpclm = -6.133346860e-08 wpclm = -4.514812308e-07 ppclm = 2.771138705e-13   pdiblc1 = 0.39   pdiblc2 = 7.442212442e-03 lpdiblc2 = 3.792036167e-09 wpdiblc2 = -7.873642851e-09 ppdiblc2 = -2.025493350e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.547765423e-03 lalpha0 = 1.311301707e-09 walpha0 = 2.193915736e-09 palpha0 = -1.045303889e-15   alpha1 = 0.0   beta0 = 1.515612294e+01 lbeta0 = 3.986444850e-06 wbeta0 = 5.398312706e-06 pbeta0 = -1.800191486e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.176829413e-01 lkt1 = -1.327937609e-08 wkt1 = -8.144748385e-08 pkt1 = 2.019475047e-14   kt2 = -1.305142721e-02 lkt2 = 3.198224575e-10 wkt2 = -5.290289901e-08 pkt2 = 8.296899551e-15   at = 6.165702106e+04 lat = -3.824167378e-04 wat = 7.457026445e-02 pat = -2.137333483e-8   ute = -1.570376333e+00 lute = -2.236563751e-07 wute = 5.155623309e-07 pute = 4.321475990e-13   ua1 = -8.110987704e-10 lua1 = -1.176222101e-16 wua1 = 4.029874337e-15 pua1 = -6.821579411e-23   ub1 = 1.566178081e-18 lub1 = -1.109181072e-25 wub1 = -5.111727976e-24 pub1 = 5.088575593e-31   uc1 = 1.001496256e-10 luc1 = -4.335963860e-17 wuc1 = -2.031314378e-16 puc1 = 8.205387908e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.46 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.244707215e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.935606067e-08 wvth0 = 7.647305581e-08 pvth0 = -2.101085689e-14   k1 = 3.970790627e-01 lk1 = 4.535967443e-08 wk1 = -2.030038938e-07 pk1 = 5.939561996e-14   k2 = -9.408034289e-03 lk2 = -1.851499056e-08 wk2 = 8.439044290e-08 pk2 = -1.842462863e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.574894221e+05 lvsat = -1.431685041e-02 wvsat = -2.661329380e-01 pvsat = 4.720578549e-8   ua = -2.405365401e-09 lua = 3.063777033e-17 wua = 4.608648823e-16 pua = -9.203032921e-23   ub = 3.163743765e-18 lub = -5.138026617e-26 wub = -1.689082559e-24 pub = 1.666925168e-31   uc = 6.866307830e-11 luc = -3.659942326e-18 wuc = 2.190121470e-18 puc = -5.291262652e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.737805106e-02 lu0 = 2.627791223e-10 wu0 = -1.477499526e-08 pu0 = 1.423941972e-15   a0 = 5.259109597e+00 la0 = -9.477178449e-07 wa0 = 2.406609183e-07 pa0 = -4.336830078e-14   keta = 1.656652093e-01 lketa = -5.152954760e-08 wketa = 3.619540325e-09 pketa = 4.214677060e-15   a1 = 0.0   a2 = 0.38689047   ags = -3.077813910e+00 lags = 7.700844294e-07 wags = 4.040491594e-07 pags = -1.010951199e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.408820716e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.815088709e-09 wvoff = -4.907484055e-08 pvoff = 1.151053979e-14   nfactor = {1.211749293e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.254274540e-07 wnfactor = -8.165123148e-07 pnfactor = 2.343421446e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.555864322e-05 lcit = 3.704770301e-12 wcit = 5.968091891e-11 pcit = -1.075479999e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.723280532e-01 leta0 = 4.670697304e-08 weta0 = -1.377019212e-08 peta0 = -1.014410158e-15   etab = -8.482788048e-02 letab = 1.368935145e-08 wetab = 1.638576489e-07 petab = -3.264076012e-14   dsub = -2.592880590e-01 ldsub = 1.064539496e-07 wdsub = 9.870193316e-07 pdsub = -1.757808175e-13   voffl = 0.0   minv = 0.0   pclm = 3.866732518e-02 lpclm = 2.443277171e-08 wpclm = 2.068283726e-06 ppclm = -3.533439205e-13   pdiblc1 = -1.163910051e+00 lpdiblc1 = 3.887960644e-07 wpdiblc1 = -2.554278431e-08 ppdiblc1 = 6.390932348e-15   pdiblc2 = 5.525877592e-02 lpdiblc2 = -8.171907097e-09 wpdiblc2 = -7.503752647e-08 ppdiblc2 = 1.477924615e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.008763796e-03 lalpha0 = -1.329994687e-09 walpha0 = -6.466729737e-09 palpha0 = 1.121632911e-15   alpha1 = 0.0   beta0 = 3.646184145e+01 lbeta0 = -1.344352450e-06 wbeta0 = -3.786633104e-06 pbeta0 = 4.979278810e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.941801173e-01 lkt1 = -1.915990018e-08 wkt1 = 1.207455154e-08 pkt1 = -3.204930398e-15   kt2 = 1.703386585e-02 lkt2 = -7.207668294e-09 wkt2 = -7.898297655e-08 pkt2 = 1.482226535e-14   at = 4.421040815e+04 lat = 3.982813045e-03 wat = -6.967226922e-02 pat = 1.471686831e-8   ute = -4.476775215e+00 lute = 5.035391572e-07 wute = 8.324106133e-06 pute = -1.521589103e-12   ua1 = -5.148021246e-09 lua1 = 9.674974779e-16 wua1 = 1.526628274e-14 pua1 = -2.879621359e-21   ub1 = 4.047525393e-18 lub1 = -7.317636113e-25 wub1 = -1.282547086e-23 pub1 = 2.438874598e-30   uc1 = -1.967170183e-10 luc1 = 3.091788004e-17 wuc1 = 3.028804865e-16 puc1 = -4.455283445e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.47 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.140718654e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.550263482e-08 wvth0 = -7.038922553e-07 pvth0 = 1.196148740e-13   k1 = 6.515973258e-01 lk1 = -5.057891655e-10 wk1 = 7.604434428e-07 pk1 = -1.142224073e-13   k2 = -1.280393624e-01 lk2 = 2.862967922e-09 wk2 = -1.880918422e-07 pk2 = 3.067804157e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.466485231e+05 lvsat = 5.657233790e-03 wvsat = -9.633702892e-04 pvsat = -5.790964571e-10   ua = -1.540135190e-09 lua = -1.252810398e-16 wua = -2.428564930e-16 pua = 3.478378121e-23   ub = 3.410055368e-18 lub = -9.576684865e-26 wub = -2.822556278e-24 pub = 3.709501483e-31   uc = 1.512507812e-10 luc = -1.854265933e-17 wuc = -1.632197271e-16 puc = 2.451641911e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.827571215e-02 lu0 = -3.503083894e-09 wu0 = -2.936499492e-08 pu0 = 4.053132862e-15   a0 = 0.0   keta = 1.582552095e-01 lketa = -5.019422859e-08 wketa = 1.622312108e-07 pketa = -2.436793902e-14   a1 = 0.0   a2 = 0.38689047   ags = 9.360418900e-01 lags = 4.676754491e-08 wags = -9.427813720e-07 pags = 1.416104760e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.733751438e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.367050279e-08 wvoff = 8.890027154e-08 pvoff = -1.335326529e-14   nfactor = {-1.402880988e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.965969038e-07 wnfactor = 6.653655243e-06 pnfactor = -1.111819400e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.003416667e-05 lcit = 4.511282004e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.255162071e-01 leta0 = -6.966051897e-09 weta0 = -1.165289209e-07 peta0 = 1.750322657e-14   etab = -5.323522497e-02 letab = 7.996196967e-09 wetab = -1.037597496e-07 petab = 1.558523319e-14   dsub = 6.891881631e-01 ldsub = -6.446620804e-08 wdsub = 6.950003742e-08 pdsub = -1.043925312e-14   voffl = 0.0   minv = 0.0   pclm = 2.054958330e-01 lpclm = -5.630559541e-09 wpclm = 6.457049439e-07 ppclm = -9.698811110e-14   pdiblc1 = 9.616217867e-01 lpdiblc1 = 5.764599521e-09 wpdiblc1 = 5.959983005e-08 ppdiblc1 = -8.952192473e-15   pdiblc2 = 3.032499028e-02 lpdiblc2 = -3.678714257e-09 wpdiblc2 = 4.190362311e-08 ppdiblc2 = -6.294133709e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.100194187e-03 lalpha0 = -2.652409002e-10 walpha0 = -1.456804030e-09 palpha0 = 2.188192493e-16   alpha1 = 0.0   beta0 = 3.420063341e+01 lbeta0 = -9.368714550e-07 wbeta0 = -6.148077918e-06 pbeta0 = 9.234720437e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.383991394e-02 lkt1 = -4.985605653e-08 wkt1 = -3.430119460e-08 pkt1 = 5.152210934e-15   kt2 = -7.960640827e-02 lkt2 = 1.020739230e-08 wkt2 = 1.963793539e-08 pkt2 = -2.949716085e-15   at = -3.770510631e+04 lat = 1.874439833e-02 wat = 7.205256783e-02 pat = -1.082265595e-8   ute = -1.778237447e+00 lute = 1.724915876e-08 wute = -7.181185769e-07 pute = 1.078650009e-13   ua1 = 5.606148783e-10 lua1 = -6.122729484e-17 wua1 = -4.285362578e-15 pua1 = 6.436828861e-22   ub1 = 3.186582166e-19 lub1 = -5.980310185e-26 wub1 = 4.255354048e-24 pub1 = -6.391754548e-31   uc1 = 4.525757967e-11 luc1 = -1.268715239e-17 wuc1 = 3.342581206e-16 puc1 = -5.020724101e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.48 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.49 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.50 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.067921137e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.801091811e-8   k1 = 6.085977213e-01 lk1 = -3.013663295e-7   k2 = -8.672152030e-02 lk2 = 1.172588584e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.584181798e+05 lvsat = -6.315050823e-1   ua = -8.491117511e-10 lua = -5.132084964e-16   ub = 2.001737703e-18 lub = 6.048601861e-25   uc = -6.766810227e-12 luc = 1.164755580e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.851148953e-02 lu0 = 4.084627936e-10   a0 = 2.012192134e+00 la0 = -3.721264076e-7   keta = 1.812485761e-01 lketa = -7.250314603e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.795138190e-01 lags = 3.349550932e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.034277124e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.722690564e-8   nfactor = {2.324936696e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.922886128e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081488e-01 leta0 = -3.180488942e-7   etab = -1.395071238e-01 letab = 2.780427440e-7   dsub = 7.177730901e-01 ldsub = -6.311247038e-7   voffl = 0.0   minv = 0.0   pclm = 1.654664607e-01 lpclm = 1.381412367e-7   pdiblc1 = 0.39   pdiblc2 = 3.389771663e-03 lpdiblc2 = 1.671817011e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.097348274e-05 lalpha0 = 3.308506342e-10 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.439514272e+01 lbeta0 = 1.359357776e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.467388838e-01 lkt1 = -4.356669758e-8   kt2 = -3.563892569e-02 lkt2 = -2.900445890e-9   at = 6.728892844e+04 lat = -3.623757086e-2   ute = -1.241906263e+00 lute = 2.444375778e-7   ua1 = 1.880891523e-09 lua1 = 3.308508622e-16   ub1 = -1.037656099e-18 lub1 = -1.713463413e-24   uc1 = 1.360335423e-10 luc1 = -2.904770555e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.51 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.311836549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.222835344e-9   k1 = 4.583800923e-01 lk1 = -9.002767689e-10   k2 = -2.395585101e-02 lk2 = -8.285347135e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.291513410e+03 lvsat = 8.282146151e-2   ua = -7.030680795e-10 lua = -8.053257785e-16   ub = 2.242211008e-18 lub = 1.238642792e-25   uc = 5.839842106e-11 luc = -1.386826347e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.361250364e-02 lu0 = -9.794611123e-9   a0 = 2.200844797e+00 la0 = -7.494704070e-7   keta = -2.499640876e-01 lketa = 1.374822657e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.122974228e+00 lags = 5.442873283e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.189297374e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.780322171e-9   nfactor = {6.288350457e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.469664874e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.500102500e-05 lcit = -1.000307521e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.665336366e-04 leta0 = -1.330809126e-10   etab = -5.280957584e-04 letab = 5.619727653e-11   dsub = 2.317195398e-01 ldsub = 3.410820376e-7   voffl = 0.0   minv = 0.0   pclm = 2.571446350e-01 lpclm = -4.523390610e-8   pdiblc1 = 0.39   pdiblc2 = 8.802396275e-03 lpdiblc2 = 5.891811299e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.018269961e-04 lalpha0 = -1.548000976e-10   alpha1 = 0.0   beta0 = 2.160961475e+01 lbeta0 = -8.368452684e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675097929e-01 lkt1 = -2.020621192e-9   kt2 = -5.146694688e-02 lkt2 = 2.875884123e-8   at = 1.978497689e+04 lat = 5.878007055e-2   ute = -1.146505494e+00 lute = 5.361648313e-8   ua1 = 2.097010394e-09 lua1 = -1.014311826e-16   ub1 = -2.063034584e-18 lub1 = 3.375037576e-25   uc1 = 3.158515721e-11 luc1 = -8.155887336e-17 wuc1 = -6.162975822e-33 puc1 = 5.877471754e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.52 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.484424942e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.039541954e-9   k1 = 4.420636819e-01 lk1 = 1.541947845e-8   k2 = -2.434789377e-02 lk2 = -7.893224012e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.699843173e+04 lvsat = 1.011151561e-1   ua = -1.165047954e-09 lua = -3.432511986e-16   ub = 2.307635860e-18 lub = 5.842601482e-26   uc = 3.230101594e-11 luc = 1.223449161e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.712875607e-02 lu0 = -3.309534390e-9   a0 = 1.925130097e+00 la0 = -4.736991857e-7   keta = -2.250661291e-01 lketa = 1.125792031e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.108400671e+00 lags = -1.441546127e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.074687619e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.683002788e-9   nfactor = {2.067502720e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.070227287e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.844132739e-03 leta0 = 2.278079649e-09 weta0 = 4.135903063e-25 peta0 = 1.972152263e-31   etab = -8.189622331e-04 letab = 3.471233788e-10   dsub = 1.452881600e-01 ldsub = 4.275311359e-7   voffl = 0.0   minv = 0.0   pclm = 9.894369870e-02 lpclm = 1.129994614e-7   pdiblc1 = 0.39   pdiblc2 = 2.204341243e-02 lpdiblc2 = -7.351919269e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.675933760e-05 lalpha0 = 9.383719628e-11 palpha0 = 1.232595164e-32   alpha1 = 0.0   beta0 = 1.726000329e+01 lbeta0 = 3.513657866e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.683795285e-01 lkt1 = -1.150707347e-9   kt2 = -9.625635970e-03 lkt2 = -1.309104714e-8   at = 7.570883437e+04 lat = 2.844748684e-3   ute = -1.056585117e+00 lute = -3.632232755e-8   ua1 = 2.530519227e-09 lua1 = -5.350288854e-16   ub1 = -2.159277735e-18 lub1 = 4.337666389e-25   uc1 = -8.822368291e-11 luc1 = 3.827452758e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.53 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.024524205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.505557715e-08 wvth0 = -2.117582368e-22   k1 = 3.451653516e-01 lk1 = 6.388850775e-8   k2 = -3.742368333e-03 lk2 = -1.820021086e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.199394048e+05 lvsat = -1.740233441e-2   ua = -1.479233181e-09 lua = -1.860941771e-16   ub = 2.549242254e-18 lub = -6.242671146e-26   uc = 7.170427229e-11 luc = -7.475214225e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.845240547e-02 lu0 = -3.971630436e-9   a0 = 4.411000044e-01 la0 = 2.686200869e-7   keta = 2.712863325e-02 lketa = -1.356987800e-8   a1 = 0.0   a2 = 0.38689047   ags = 4.531657218e-01 lags = -1.133843294e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.340416673e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.608897350e-9   nfactor = {1.667665112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.307030435e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.100000000e-09 lcit = 2.503075841e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.551186649e-03 leta0 = 7.951891478e-11   etab = 8.363960144e-03 letab = -4.246220309e-09 wetab = 1.344168495e-24 petab = 5.669937756e-31   dsub = 1.651174065e+00 ldsub = -3.257205233e-7   voffl = 0.0   minv = 0.0   pclm = 9.072817740e-02 lpclm = 1.171089063e-7   pdiblc1 = 0.39   pdiblc2 = 2.372125092e-03 lpdiblc2 = 2.487757016e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.135033778e-03 lalpha0 = 6.381975126e-10 walpha0 = 1.033975766e-25 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.863226702e+01 lbeta0 = 2.827244687e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.701295490e-01 lkt1 = -2.753383425e-10   kt2 = -4.711727502e-02 lkt2 = 5.662458166e-9   at = 1.096751699e+05 lat = -1.414538219e-2   ute = -1.238389462e+00 lute = 5.461711484e-8   ua1 = 1.783864614e-09 lua1 = -1.615485147e-16   ub1 = -1.725425035e-18 lub1 = 2.167513493e-25   uc1 = -3.065312391e-11 luc1 = 9.477446116e-18 wuc1 = -6.162975822e-33   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.54 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.737141378e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.288561513e-8   k1 = 2.663584429e-01 lk1 = 8.360639035e-8   k2 = 4.493363768e-02 lk2 = -3.037919095e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.611801649e+04 lvsat = 1.608044604e-2   ua = -2.108599945e-09 lua = -2.862346577e-17   ub = 2.076090149e-18 lub = 5.595831101e-26   uc = 7.007336669e-11 luc = -7.067153491e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.863964893e-03 lu0 = 1.179700338e-9   a0 = 5.414078764e+00 la0 = -9.756440637e-7   keta = 1.679959457e-01 lketa = -4.881558391e-08 pketa = 6.310887242e-30   a1 = 0.0   a2 = 0.38689047   ags = -2.817633893e+00 lags = 7.049860882e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.724829116e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.522708888e-8   nfactor = {6.859712211e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.763277635e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.287178571e-05 lcit = -3.220585145e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.811951149e-01 leta0 = 4.605376229e-08 weta0 = 2.316105715e-23 peta0 = -3.155443621e-30   etab = 2.068523573e-02 letab = -7.329065066e-09 petab = -1.577721810e-30   dsub = 3.762848673e-01 ldsub = -6.736871535e-9   voffl = 0.0   minv = 0.0   pclm = 1.370500551e+00 lpclm = -2.030965404e-7   pdiblc1 = -1.180357857e+00 lpdiblc1 = 3.929113876e-7   pdiblc2 = 6.939742286e-03 lpdiblc2 = 1.344916356e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.844632243e-03 lalpha0 = -6.077398241e-10   alpha1 = 0.0   beta0 = 3.402350878e+01 lbeta0 = -1.023720959e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.864049321e-01 lkt1 = -2.122365610e-8   kt2 = -3.382576771e-02 lkt2 = 2.336856581e-9   at = -6.537668571e+02 lat = 1.345946944e-2   ute = 8.833796714e-01 lute = -4.762601312e-7   ua1 = 4.682420453e-09 lua1 = -8.867816784e-16 pua1 = 1.880790961e-37   ub1 = -4.211200436e-18 lub1 = 8.387047834e-25   uc1 = -1.682705457e-12 luc1 = 2.228902567e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.55 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.781151963e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.827921335e-10 wvth0 = -1.821649863e-07 pvth0 = 3.282704136e-14   k1 = 1.241219099e+00 lk1 = -9.206837413e-08 wk1 = -1.552155857e-07 pk1 = 2.797062462e-14   k2 = -2.895536230e-01 lk2 = 2.989708587e-08 wk2 = 6.273334394e-08 pk2 = -1.130486225e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.298987478e+05 lvsat = 8.190939348e-03 wvsat = 2.504836070e-02 pvsat = -4.513839840e-9   ua = 1.972315546e-10 lua = -4.441458311e-16 wua = -2.940917553e-15 pua = 5.299680476e-22   ub = 6.872292308e-19 lub = 3.062379927e-25 wub = 1.405883800e-24 pub = -2.533472902e-31   uc = -8.001211550e-11 luc = 1.997900083e-17 wuc = 1.959223010e-16 puc = -3.530617825e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 5.199346314e-02 lu0 = -6.772655893e-09 wu0 = -5.066811350e-08 pu0 = 9.130647394e-15   a0 = 0.0   keta = 1.486278340e+00 lketa = -2.863766629e-07 wketa = -1.900135591e-06 pketa = 3.424139341e-13   a1 = 0.0   a2 = 0.38689047   ags = 3.178266412e-01 lags = 1.399604226e-07 wags = 1.728218073e-08 pags = -3.114335379e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-3.286547524e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.337003545e-08 wvoff = 3.300432926e-07 pvoff = -5.947545154e-14   nfactor = {3.327217149e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.620411135e-10 wnfactor = -6.919979590e-07 pnfactor = 1.247014922e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.003416667e-05 lcit = 4.511282004e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.659846883e-01 leta0 = 4.331276737e-08 weta0 = 3.361603096e-07 peta0 = -6.057776860e-14   etab = -2.013226437e-01 letab = 3.267786485e-08 wetab = 1.262140882e-07 petab = -2.274440976e-14   dsub = 7.339414326e-01 ldsub = -7.118837288e-8   voffl = 0.0   minv = 0.0   pclm = 1.750484899e+00 lpclm = -2.715716199e-07 wpclm = -1.753601276e-06 ppclm = 3.160077180e-13   pdiblc1 = 6.520971522e-01 lpdiblc1 = 6.269383269e-08 wpdiblc1 = 5.402792066e-07 ppdiblc1 = -9.736101442e-14   pdiblc2 = 6.916690955e-02 lpdiblc2 = -9.868730321e-09 wpdiblc2 = -1.841632384e-08 ppdiblc2 = 3.318713638e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.289096887e-04 lalpha0 = 6.185195881e-11 walpha0 = 1.604521945e-09 palpha0 = -2.891428771e-16   alpha1 = 0.0   beta0 = 2.274853840e+01 lbeta0 = 1.008085079e-06 wbeta0 = 1.163656755e-05 pbeta0 = -2.096967655e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 3.899635466e-01 lkt1 = -1.250881378e-07 wkt1 = -6.769214166e-07 pkt1 = 1.219846239e-13   kt2 = -4.105158873e-02 lkt2 = 3.638985657e-09 wkt2 = -4.023615716e-08 pkt2 = 7.250756701e-15   at = -8.379332199e+04 lat = 2.844163297e-02 wat = 1.436257233e-01 pat = -2.588207346e-8   ute = -2.177363100e+00 lute = 7.530101996e-08 wute = -9.829240292e-08 pute = 1.771278247e-14   ua1 = -4.034935794e-09 lua1 = 6.841295041e-16 wua1 = 2.851343794e-15 pua1 = -5.138264084e-22   ub1 = 6.218729861e-18 lub1 = -1.040820806e-24 wub1 = -4.907221213e-24 pub1 = 8.843057986e-31   uc1 = 4.420312853e-10 luc1 = -7.773057713e-17 wuc1 = -2.819155732e-16 puc1 = 5.080259587e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.56 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.57 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.58 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.067921137e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.801091811e-8   k1 = 6.085977213e-01 lk1 = -3.013663295e-7   k2 = -8.672152030e-02 lk2 = 1.172588584e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.584181798e+05 lvsat = -6.315050823e-1   ua = -8.491117511e-10 lua = -5.132084964e-16   ub = 2.001737703e-18 lub = 6.048601861e-25   uc = -6.766810227e-12 luc = 1.164755580e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.851148953e-02 lu0 = 4.084627936e-10   a0 = 2.012192134e+00 la0 = -3.721264076e-7   keta = 1.812485761e-01 lketa = -7.250314603e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.795138190e-01 lags = 3.349550932e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.034277124e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.722690564e-8   nfactor = {2.324936696e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.922886128e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081488e-01 leta0 = -3.180488942e-7   etab = -1.395071238e-01 letab = 2.780427440e-7   dsub = 7.177730901e-01 ldsub = -6.311247038e-7   voffl = 0.0   minv = 0.0   pclm = 1.654664607e-01 lpclm = 1.381412367e-7   pdiblc1 = 0.39   pdiblc2 = 3.389771663e-03 lpdiblc2 = 1.671817011e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.097348274e-05 lalpha0 = 3.308506342e-10 palpha0 = 9.860761315e-32   alpha1 = 0.0   beta0 = 1.439514272e+01 lbeta0 = 1.359357776e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.467388838e-01 lkt1 = -4.356669758e-8   kt2 = -3.563892569e-02 lkt2 = -2.900445890e-9   at = 6.728892845e+04 lat = -3.623757086e-2   ute = -1.241906263e+00 lute = 2.444375778e-7   ua1 = 1.880891523e-09 lua1 = 3.308508622e-16   ub1 = -1.037656099e-18 lub1 = -1.713463413e-24   uc1 = 1.360335423e-10 luc1 = -2.904770555e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.59 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.311836549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.222835344e-9   k1 = 4.583800923e-01 lk1 = -9.002767689e-10   k2 = -2.395585101e-02 lk2 = -8.285347135e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.291513410e+03 lvsat = 8.282146151e-2   ua = -7.030680795e-10 lua = -8.053257785e-16   ub = 2.242211008e-18 lub = 1.238642792e-25   uc = 5.839842106e-11 luc = -1.386826347e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.361250364e-02 lu0 = -9.794611123e-9   a0 = 2.200844797e+00 la0 = -7.494704070e-7   keta = -2.499640876e-01 lketa = 1.374822657e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.122974228e+00 lags = 5.442873283e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.189297374e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.780322171e-9   nfactor = {6.288350457e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.469664874e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.500102500e-05 lcit = -1.000307521e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.665336366e-04 leta0 = -1.330809126e-10   etab = -5.280957584e-04 letab = 5.619727653e-11   dsub = 2.317195398e-01 ldsub = 3.410820376e-7   voffl = 0.0   minv = 0.0   pclm = 2.571446350e-01 lpclm = -4.523390610e-8   pdiblc1 = 0.39   pdiblc2 = 8.802396275e-03 lpdiblc2 = 5.891811299e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.018269961e-04 lalpha0 = -1.548000976e-10   alpha1 = 0.0   beta0 = 2.160961475e+01 lbeta0 = -8.368452684e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675097929e-01 lkt1 = -2.020621192e-9   kt2 = -5.146694687e-02 lkt2 = 2.875884123e-8   at = 1.978497689e+04 lat = 5.878007055e-2   ute = -1.146505494e+00 lute = 5.361648313e-8   ua1 = 2.097010394e-09 lua1 = -1.014311826e-16   ub1 = -2.063034584e-18 lub1 = 3.375037576e-25   uc1 = 3.158515721e-11 luc1 = -8.155887336e-17 puc1 = 1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.60 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.484424942e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.039541954e-9   k1 = 4.420636819e-01 lk1 = 1.541947845e-8   k2 = -2.434789377e-02 lk2 = -7.893224012e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.699843173e+04 lvsat = 1.011151561e-1   ua = -1.165047954e-09 lua = -3.432511986e-16   ub = 2.307635860e-18 lub = 5.842601482e-26   uc = 3.230101594e-11 luc = 1.223449161e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.712875607e-02 lu0 = -3.309534390e-9   a0 = 1.925130097e+00 la0 = -4.736991857e-7   keta = -2.250661291e-01 lketa = 1.125792031e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.108400671e+00 lags = -1.441546127e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.074687619e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.683002788e-9   nfactor = {2.067502720e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.070227287e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.844132739e-03 leta0 = 2.278079649e-09 peta0 = 7.888609052e-31   etab = -8.189622331e-04 letab = 3.471233788e-10   dsub = 1.452881600e-01 ldsub = 4.275311359e-7   voffl = 0.0   minv = 0.0   pclm = 9.894369870e-02 lpclm = 1.129994614e-7   pdiblc1 = 0.39   pdiblc2 = 2.204341243e-02 lpdiblc2 = -7.351919269e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.675933760e-05 lalpha0 = 9.383719628e-11 palpha0 = 2.465190329e-32   alpha1 = 0.0   beta0 = 1.726000329e+01 lbeta0 = 3.513657866e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.683795285e-01 lkt1 = -1.150707347e-9   kt2 = -9.625635970e-03 lkt2 = -1.309104714e-8   at = 7.570883437e+04 lat = 2.844748684e-3   ute = -1.056585117e+00 lute = -3.632232755e-8   ua1 = 2.530519227e-09 lua1 = -5.350288854e-16   ub1 = -2.159277735e-18 lub1 = 4.337666389e-25   uc1 = -8.822368291e-11 luc1 = 3.827452758e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.61 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.024524205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.505557715e-08 wvth0 = 4.235164736e-22   k1 = 3.451653516e-01 lk1 = 6.388850775e-8   k2 = -3.742368333e-03 lk2 = -1.820021086e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.199394048e+05 lvsat = -1.740233441e-2   ua = -1.479233181e-09 lua = -1.860941771e-16   ub = 2.549242254e-18 lub = -6.242671146e-26   uc = 7.170427229e-11 luc = -7.475214225e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.845240547e-02 lu0 = -3.971630436e-9   a0 = 4.411000044e-01 la0 = 2.686200869e-7   keta = 2.712863325e-02 lketa = -1.356987800e-8   a1 = 0.0   a2 = 0.38689047   ags = 4.531657218e-01 lags = -1.133843294e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.340416673e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.608897350e-9   nfactor = {1.667665112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.307030435e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.100000000e-09 lcit = 2.503075841e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.551186649e-03 leta0 = 7.951891478e-11   etab = 8.363960144e-03 letab = -4.246220309e-09 wetab = 1.033975766e-24 petab = 5.916456789e-31   dsub = 1.651174065e+00 ldsub = -3.257205233e-7   voffl = 0.0   minv = 0.0   pclm = 9.072817740e-02 lpclm = 1.171089063e-7   pdiblc1 = 0.39   pdiblc2 = 2.372125092e-03 lpdiblc2 = 2.487757016e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.135033778e-03 lalpha0 = 6.381975126e-10 walpha0 = 4.135903063e-25 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.863226702e+01 lbeta0 = 2.827244687e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.701295490e-01 lkt1 = -2.753383425e-10   kt2 = -4.711727502e-02 lkt2 = 5.662458166e-9   at = 1.096751699e+05 lat = -1.414538219e-2   ute = -1.238389462e+00 lute = 5.461711484e-8   ua1 = 1.783864614e-09 lua1 = -1.615485147e-16   ub1 = -1.725425035e-18 lub1 = 2.167513493e-25   uc1 = -3.065312391e-11 luc1 = 9.477446116e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.62 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.737141378e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.288561513e-8   k1 = 2.663584429e-01 lk1 = 8.360639035e-8   k2 = 4.493363768e-02 lk2 = -3.037919095e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.611801649e+04 lvsat = 1.608044604e-2   ua = -2.108599945e-09 lua = -2.862346577e-17   ub = 2.076090149e-18 lub = 5.595831101e-26   uc = 7.007336669e-11 luc = -7.067153491e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.863964893e-03 lu0 = 1.179700338e-9   a0 = 5.414078764e+00 la0 = -9.756440637e-7   keta = 1.679959457e-01 lketa = -4.881558391e-08 wketa = -5.293955920e-23   a1 = 0.0   a2 = 0.38689047   ags = -2.817633893e+00 lags = 7.049860882e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.724829116e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.522708888e-8   nfactor = {6.859712211e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.763277635e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.287178571e-05 lcit = -3.220585145e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.811951149e-01 leta0 = 4.605376229e-08 weta0 = 2.646977960e-23 peta0 = 1.262177448e-29   etab = 2.068523573e-02 letab = -7.329065066e-9   dsub = 3.762848673e-01 ldsub = -6.736871535e-9   voffl = 0.0   minv = 0.0   pclm = 1.370500551e+00 lpclm = -2.030965404e-7   pdiblc1 = -1.180357857e+00 lpdiblc1 = 3.929113876e-7   pdiblc2 = 6.939742286e-03 lpdiblc2 = 1.344916356e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.844632243e-03 lalpha0 = -6.077398241e-10   alpha1 = 0.0   beta0 = 3.402350878e+01 lbeta0 = -1.023720959e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.864049321e-01 lkt1 = -2.122365610e-8   kt2 = -3.382576771e-02 lkt2 = 2.336856581e-9   at = -6.537668571e+02 lat = 1.345946944e-2   ute = 8.833796714e-01 lute = -4.762601312e-7   ua1 = 4.682420453e-09 lua1 = -8.867816784e-16   ub1 = -4.211200436e-18 lub1 = 8.387047834e-25 pub1 = -3.503246161e-46   uc1 = -1.682705457e-12 luc1 = 2.228902567e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.63 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-7.593204303e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.873338792e-07 wvth0 = 7.545978870e-07 pvth0 = -1.359823122e-13   k1 = 2.359654982e+00 lk1 = -2.936161125e-07 wk1 = -1.165118451e-06 pk1 = 2.099601705e-13   k2 = -2.824602511e-01 lk2 = 2.861882478e-08 wk2 = 5.632831281e-08 pk2 = -1.015064361e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.336389603e+05 lvsat = 5.568175205e-02 wvsat = 2.630123697e-01 pvsat = -4.739614408e-8   ua = -8.185212132e-09 lua = 1.066412433e-15 wua = 4.628093799e-15 pua = -8.340056430e-22   ub = 2.161201879e-18 lub = 4.062075159e-26 wub = 7.494545713e-26 pub = -1.350554610e-32   uc = 2.537635184e-11 luc = 9.874720697e-19 wuc = 1.007607305e-16 puc = -1.815758745e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.282335827e-01 lu0 = 2.570515890e-08 wu0 = 1.120696998e-07 pu0 = -2.019552026e-14   a0 = 0.0   keta = -3.124562033e+00 lketa = 5.445198266e-07 wketa = 2.263268833e-06 pketa = -4.078523600e-13   a1 = 0.0   a2 = 0.38689047   ags = 2.741931941e-01 lags = 1.478233880e-07 wags = 5.668143817e-08 pags = -1.021427857e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {7.417219217e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.495171931e-07 wvoff = -6.364640291e-07 pvoff = 1.146940004e-13   nfactor = {1.399650819e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.922297551e-06 wnfactor = -1.032594100e-05 pnfactor = 1.860786198e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.003416667e-05 lcit = 4.511282004e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.317879176e-01 leta0 = 5.517083830e-08 weta0 = 3.955779936e-07 peta0 = -7.128513233e-14   etab = 1.619018962e-01 letab = -3.277701336e-08 wetab = -2.017631423e-07 petab = 3.635872707e-14   dsub = 7.348430378e-01 ldsub = -7.135084664e-08 wdsub = -8.141133971e-10 pdsub = 1.467073047e-16   voffl = 0.0   minv = 0.0   pclm = -1.999434713e-01 lpclm = 7.990532460e-08 wpclm = 7.557525089e-09 ppclm = -1.361903809e-15   pdiblc1 = 2.413355319e+00 lpdiblc1 = -2.546936953e-07 wpdiblc1 = -1.050066468e-06 ppdiblc1 = 1.892272279e-13   pdiblc2 = 3.094720034e-01 lpdiblc2 = -5.317290975e-08 wpdiblc2 = -2.354022113e-07 ppdiblc2 = 4.242065549e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.236432901e-03 lalpha0 = 4.880985202e-10 walpha0 = 3.740331690e-09 palpha0 = -6.740264722e-16   alpha1 = 0.0   beta0 = -1.105095479e+02 lbeta0 = 2.502185852e-05 wbeta0 = 1.319632891e-04 pbeta0 = -2.378044452e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -9.223371618e-01 lkt1 = 1.113950113e-07 wkt1 = 5.080336310e-07 pkt1 = -9.155020047e-14   kt2 = -3.545148020e-01 lkt2 = 6.012662401e-08 wkt2 = 2.428085859e-07 pkt2 = -4.375532123e-14   at = 1.606388557e+05 lat = -1.560626761e-02 wat = -7.708675591e-02 pat = 1.389141885e-8   ute = -3.906690238e+00 lute = 3.869344169e-07 wute = 1.463220830e-06 pute = -2.636797096e-13   ua1 = -3.580582124e-09 lua1 = 6.022527009e-16 wua1 = 2.441080604e-15 pua1 = -4.398949302e-22   ub1 = 1.657060898e-19 lub1 = 4.996434293e-26 wub1 = 5.584171316e-25 pub1 = -1.006295592e-31   uc1 = 8.766536264e-10 luc1 = -1.560516961e-16 wuc1 = -6.743621623e-16 puc1 = 1.215234335e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.64 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.65 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.66 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.067921137e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.801091811e-8   k1 = 6.085977213e-01 lk1 = -3.013663295e-7   k2 = -8.672152030e-02 lk2 = 1.172588584e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.584181798e+05 lvsat = -6.315050823e-1   ua = -8.491117511e-10 lua = -5.132084964e-16   ub = 2.001737703e-18 lub = 6.048601861e-25   uc = -6.766810227e-12 luc = 1.164755580e-16 puc = 2.350988702e-38   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.851148953e-02 lu0 = 4.084627936e-10   a0 = 2.012192134e+00 la0 = -3.721264076e-7   keta = 1.812485761e-01 lketa = -7.250314603e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.795138190e-01 lags = 3.349550932e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.034277124e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.722690564e-8   nfactor = {2.324936696e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.922886128e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081488e-01 leta0 = -3.180488942e-7   etab = -1.395071238e-01 letab = 2.780427440e-7   dsub = 7.177730901e-01 ldsub = -6.311247038e-7   voffl = 0.0   minv = 0.0   pclm = 1.654664607e-01 lpclm = 1.381412367e-7   pdiblc1 = 0.39   pdiblc2 = 3.389771663e-03 lpdiblc2 = 1.671817011e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.097348274e-05 lalpha0 = 3.308506342e-10 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.439514272e+01 lbeta0 = 1.359357776e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.467388838e-01 lkt1 = -4.356669758e-8   kt2 = -3.563892569e-02 lkt2 = -2.900445890e-9   at = 6.728892845e+04 lat = -3.623757086e-2   ute = -1.241906263e+00 lute = 2.444375778e-7   ua1 = 1.880891523e-09 lua1 = 3.308508622e-16   ub1 = -1.037656099e-18 lub1 = -1.713463413e-24   uc1 = 1.360335423e-10 luc1 = -2.904770555e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.67 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.311836549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.222835344e-9   k1 = 4.583800923e-01 lk1 = -9.002767689e-10   k2 = -2.395585101e-02 lk2 = -8.285347135e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.291513410e+03 lvsat = 8.282146151e-2   ua = -7.030680795e-10 lua = -8.053257785e-16   ub = 2.242211008e-18 lub = 1.238642792e-25   uc = 5.839842106e-11 luc = -1.386826347e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.361250364e-02 lu0 = -9.794611123e-9   a0 = 2.200844797e+00 la0 = -7.494704070e-7   keta = -2.499640876e-01 lketa = 1.374822657e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.122974228e+00 lags = 5.442873283e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.189297374e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.780322171e-9   nfactor = {6.288350457e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.469664874e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.500102500e-05 lcit = -1.000307521e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.665336366e-04 leta0 = -1.330809126e-10   etab = -5.280957584e-04 letab = 5.619727653e-11   dsub = 2.317195398e-01 ldsub = 3.410820376e-7   voffl = 0.0   minv = 0.0   pclm = 2.571446350e-01 lpclm = -4.523390610e-8   pdiblc1 = 0.39   pdiblc2 = 8.802396275e-03 lpdiblc2 = 5.891811299e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.018269961e-04 lalpha0 = -1.548000976e-10   alpha1 = 0.0   beta0 = 2.160961475e+01 lbeta0 = -8.368452684e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675097930e-01 lkt1 = -2.020621192e-9   kt2 = -5.146694688e-02 lkt2 = 2.875884123e-8   at = 1.978497689e+04 lat = 5.878007055e-2   ute = -1.146505494e+00 lute = 5.361648313e-8   ua1 = 2.097010394e-09 lua1 = -1.014311826e-16   ub1 = -2.063034584e-18 lub1 = 3.375037576e-25   uc1 = 3.158515721e-11 luc1 = -8.155887336e-17 wuc1 = 6.162975822e-33 puc1 = -1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.68 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.484424942e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.039541954e-9   k1 = 4.420636819e-01 lk1 = 1.541947845e-8   k2 = -2.434789377e-02 lk2 = -7.893224012e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.699843173e+04 lvsat = 1.011151561e-1   ua = -1.165047954e-09 lua = -3.432511986e-16   ub = 2.307635860e-18 lub = 5.842601482e-26   uc = 3.230101594e-11 luc = 1.223449161e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.712875608e-02 lu0 = -3.309534390e-9   a0 = 1.925130097e+00 la0 = -4.736991857e-7   keta = -2.250661291e-01 lketa = 1.125792031e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.108400671e+00 lags = -1.441546127e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.074687619e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.683002788e-9   nfactor = {2.067502720e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.070227287e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.844132739e-03 leta0 = 2.278079649e-09 weta0 = 2.067951531e-25 peta0 = -1.972152263e-31   etab = -8.189622331e-04 letab = 3.471233788e-10   dsub = 1.452881600e-01 ldsub = 4.275311359e-7   voffl = 0.0   minv = 0.0   pclm = 9.894369870e-02 lpclm = 1.129994614e-7   pdiblc1 = 0.39   pdiblc2 = 2.204341243e-02 lpdiblc2 = -7.351919269e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.675933760e-05 lalpha0 = 9.383719628e-11   alpha1 = 0.0   beta0 = 1.726000329e+01 lbeta0 = 3.513657866e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.683795285e-01 lkt1 = -1.150707347e-9   kt2 = -9.625635970e-03 lkt2 = -1.309104714e-8   at = 7.570883437e+04 lat = 2.844748684e-3   ute = -1.056585117e+00 lute = -3.632232755e-8   ua1 = 2.530519227e-09 lua1 = -5.350288854e-16   ub1 = -2.159277735e-18 lub1 = 4.337666389e-25   uc1 = -8.822368291e-11 luc1 = 3.827452758e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.69 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.024524205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.505557715e-8   k1 = 3.451653516e-01 lk1 = 6.388850775e-8   k2 = -3.742368333e-03 lk2 = -1.820021086e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.199394048e+05 lvsat = -1.740233441e-2   ua = -1.479233181e-09 lua = -1.860941771e-16   ub = 2.549242254e-18 lub = -6.242671146e-26   uc = 7.170427229e-11 luc = -7.475214225e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.845240547e-02 lu0 = -3.971630436e-9   a0 = 4.411000044e-01 la0 = 2.686200869e-7   keta = 2.712863325e-02 lketa = -1.356987800e-8   a1 = 0.0   a2 = 0.38689047   ags = 4.531657218e-01 lags = -1.133843294e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.340416673e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.608897350e-9   nfactor = {1.667665112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.307030435e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.100000000e-09 lcit = 2.503075840e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.551186649e-03 leta0 = 7.951891478e-11   etab = 8.363960144e-03 letab = -4.246220309e-09 wetab = 1.447566072e-24 petab = 6.162975822e-31   dsub = 1.651174065e+00 ldsub = -3.257205233e-7   voffl = 0.0   minv = 0.0   pclm = 9.072817740e-02 lpclm = 1.171089063e-7   pdiblc1 = 0.39   pdiblc2 = 2.372125092e-03 lpdiblc2 = 2.487757016e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.135033778e-03 lalpha0 = 6.381975126e-10   alpha1 = 0.0   beta0 = 1.863226702e+01 lbeta0 = 2.827244687e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.701295490e-01 lkt1 = -2.753383425e-10   kt2 = -4.711727502e-02 lkt2 = 5.662458166e-9   at = 1.096751699e+05 lat = -1.414538219e-2   ute = -1.238389462e+00 lute = 5.461711484e-8   ua1 = 1.783864614e-09 lua1 = -1.615485147e-16 wua1 = -7.888609052e-31   ub1 = -1.725425035e-18 lub1 = 2.167513493e-25   uc1 = -3.065312391e-11 luc1 = 9.477446116e-18 puc1 = 1.469367939e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.70 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.737141378e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.288561513e-8   k1 = 2.663584429e-01 lk1 = 8.360639035e-8   k2 = 4.493363768e-02 lk2 = -3.037919095e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.611801649e+04 lvsat = 1.608044604e-2   ua = -2.108599945e-09 lua = -2.862346577e-17   ub = 2.076090149e-18 lub = 5.595831101e-26   uc = 7.007336669e-11 luc = -7.067153491e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.863964893e-03 lu0 = 1.179700338e-9   a0 = 5.414078764e+00 la0 = -9.756440637e-7   keta = 1.679959457e-01 lketa = -4.881558391e-08 wketa = 2.646977960e-23 pketa = -6.310887242e-30   a1 = 0.0   a2 = 0.38689047   ags = -2.817633893e+00 lags = 7.049860882e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.724829116e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.522708888e-8   nfactor = {6.859712211e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.763277635e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.287178571e-05 lcit = -3.220585145e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.811951149e-01 leta0 = 4.605376229e-08 weta0 = 3.308722450e-24 peta0 = -4.733165431e-30   etab = 2.068523573e-02 letab = -7.329065066e-09 petab = 1.577721810e-30   dsub = 3.762848673e-01 ldsub = -6.736871535e-9   voffl = 0.0   minv = 0.0   pclm = 1.370500551e+00 lpclm = -2.030965404e-7   pdiblc1 = -1.180357857e+00 lpdiblc1 = 3.929113876e-7   pdiblc2 = 6.939742286e-03 lpdiblc2 = 1.344916356e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.844632243e-03 lalpha0 = -6.077398241e-10   alpha1 = 0.0   beta0 = 3.402350878e+01 lbeta0 = -1.023720959e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.864049321e-01 lkt1 = -2.122365610e-8   kt2 = -3.382576771e-02 lkt2 = 2.336856581e-9   at = -6.537668571e+02 lat = 1.345946944e-2   ute = 8.833796714e-01 lute = -4.762601312e-7   ua1 = 4.682420453e-09 lua1 = -8.867816784e-16   ub1 = -4.211200436e-18 lub1 = 8.387047834e-25 pub1 = -1.751623080e-46   uc1 = -1.682705457e-12 luc1 = 2.228902567e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.71 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.347588160e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 8.195828634e-09 wvth0 = 1.603677020e-08 pvth0 = -2.889906174e-15   k1 = 7.914434350e-01 lk1 = -1.101655065e-8   k2 = -1.966128710e-01 lk2 = 1.314869766e-08 wk2 = -7.452856681e-09 pk2 = 1.343042038e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.970056188e+05 lvsat = -3.902054338e-03 wvsat = 1.735667314e-02 pvsat = -3.127759283e-9   ua = -1.977125981e-09 lua = -5.231573153e-17 wua = 1.573411151e-17 pua = -2.835365565e-24   ub = -1.141407489e-20 lub = 4.321370096e-25 wub = 1.689112207e-24 pub = -3.043864652e-31   uc = 1.609970186e-10 luc = -2.345205018e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.432664749e-02 lu0 = 1.509262026e-11 wu0 = 6.153151187e-09 pu0 = -1.108828610e-15   a0 = 0.0   keta = 5.301539918e-01 lketa = -1.140782746e-07 wketa = -4.520389848e-07 pketa = 8.145968525e-14   a1 = 0.0   a2 = 0.38689047   ags = 3.504845667e-01 lags = 1.340753012e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.149404927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.857657292e-09 wvoff = 1.878362253e-12 pvoff = -3.384902698e-19   nfactor = {1.373598020e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.524139762e-07 wnfactor = -9.476236579e-07 pnfactor = 1.707665213e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.003416667e-05 lcit = 4.511282004e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.006471981e-01 leta0 = -4.077663172e-8   etab = -1.096647324e-01 letab = 1.616065094e-8   dsub = 7.337472676e-01 ldsub = -7.115338338e-8   voffl = 0.0   minv = 0.0   pclm = -4.124172759e-01 lpclm = 1.181941666e-07 wpclm = 1.654170629e-07 ppclm = -2.980898182e-14   pdiblc1 = 1.0   pdiblc2 = -1.692728161e-02 lpdiblc2 = 5.645873398e-09 wpdiblc2 = 7.099401418e-09 ppdiblc2 = -1.279347633e-15   pdiblcb = 0.0   drout = -2.975549858e+01 ldrout = 5.991834015e-06 wdrout = 2.470349324e-05 pdrout = -4.451693000e-12   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.763419077e-03 lalpha0 = -4.128998054e-10 walpha0 = 2.564166450e-11 palpha0 = -4.620756151e-18   alpha1 = 0.0   beta0 = 5.918429073e+01 lbeta0 = -5.557819670e-06 wbeta0 = 5.887554804e-06 pbeta0 = -1.060966813e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.288361309e-01 lkt1 = 2.246365806e-08 wkt1 = 1.413821051e-07 pkt1 = -2.547776224e-14   kt2 = -2.770234117e-02 lkt2 = 1.233384500e-9   at = 1.185655860e+05 lat = -8.024454053e-03 wat = -4.582799948e-02 pat = 8.258434647e-9   ute = -1.937242583e+00 lute = 3.203010223e-8   ua1 = -2.949670117e-10 lua1 = 1.016842964e-17   ub1 = 9.173173900e-19 lub1 = -8.547977141e-26   uc1 = -3.101591483e-11 luc1 = 7.514893563e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.72 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.73 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4212941+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.057408308   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.774073e-10   ub = 2.152945e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.0286136   a0 = 1.9191653   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.557831   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.8442398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.74 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.067921137e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.801091811e-8   k1 = 6.085977213e-01 lk1 = -3.013663295e-7   k2 = -8.672152030e-02 lk2 = 1.172588584e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.584181798e+05 lvsat = -6.315050823e-1   ua = -8.491117511e-10 lua = -5.132084964e-16   ub = 2.001737703e-18 lub = 6.048601861e-25   uc = -6.766810227e-12 luc = 1.164755580e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.851148953e-02 lu0 = 4.084627936e-10   a0 = 2.012192134e+00 la0 = -3.721264076e-7   keta = 1.812485761e-01 lketa = -7.250314603e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.795138190e-01 lags = 3.349550932e-06 pags = -8.077935669e-28   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.034277124e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.722690564e-8   nfactor = {2.324936696e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.922886128e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.595081488e-01 leta0 = -3.180488942e-7   etab = -1.395071238e-01 letab = 2.780427440e-7   dsub = 7.177730901e-01 ldsub = -6.311247038e-7   voffl = 0.0   minv = 0.0   pclm = 1.654664607e-01 lpclm = 1.381412367e-7   pdiblc1 = 0.39   pdiblc2 = 3.389771663e-03 lpdiblc2 = 1.671817011e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.097348274e-05 lalpha0 = 3.308506342e-10   alpha1 = 0.0   beta0 = 1.439514272e+01 lbeta0 = 1.359357776e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.467388838e-01 lkt1 = -4.356669758e-8   kt2 = -3.563892569e-02 lkt2 = -2.900445890e-9   at = 6.728892844e+04 lat = -3.623757086e-2   ute = -1.241906263e+00 lute = 2.444375778e-7   ua1 = 1.880891523e-09 lua1 = 3.308508622e-16   ub1 = -1.037656099e-18 lub1 = -1.713463413e-24   uc1 = 1.360335423e-10 luc1 = -2.904770555e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.75 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.135122365e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.445897950e-07 wvth0 = 6.389087339e-08 pvth0 = -1.277948444e-13   k1 = 5.701834695e-01 lk1 = -2.245299509e-07 wk1 = -6.070476169e-08 pk1 = 1.214219679e-13   k2 = -7.548104902e-02 lk2 = 9.477561155e-08 wk2 = 2.797612151e-08 pk2 = -5.595797813e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.937312298e+04 lvsat = 6.650435631e-03 wvsat = -2.067679073e-02 pvsat = 4.135782021e-8   ua = 9.348211932e-10 lua = -4.081440091e-15 wua = -8.893083595e-16 pua = 1.778799027e-21   ub = 5.028912547e-19 lub = 3.602860346e-24 wub = 9.443810531e-25 pub = -1.888955704e-30   uc = -3.896767179e-11 luc = 1.808838823e-16 wuc = 5.286589377e-17 puc = -1.057426251e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.655545031e-02 lu0 = 4.320942239e-09 wu0 = 3.831697678e-09 pu0 = -7.664180853e-15   a0 = 2.745877452e+00 la0 = -1.839647448e-06 wa0 = -2.959309301e-07 pa0 = 5.919225261e-13   keta = -3.380073594e-01 lketa = 3.135868582e-07 wketa = 4.780397488e-08 pketa = -9.561774957e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.583829661e+00 lags = -3.775180146e-07 wags = -2.502260663e-07 pags = 5.005034290e-13   b0 = 5.712996524e-07 lb0 = -1.142716421e-12 wb0 = -3.101928593e-13 pb0 = 6.204493081e-19   b1 = 2.176415585e-07 lb1 = -4.353277335e-13 wb1 = -1.181706606e-13 pb1 = 2.363655462e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.944721734e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.548806805e-07 wvoff = 4.101652108e-08 pvoff = -8.204145055e-14   nfactor = {-1.264731687e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.257186521e-06 wnfactor = 1.028130993e-06 pnfactor = -2.056472753e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 4.017062816e-05 lcit = -6.034744129e-11 wcit = -1.366608773e-11 pcit = 2.733497701e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.292654338e-03 leta0 = 3.585676170e-09 weta0 = 1.009464703e-09 peta0 = -2.019136346e-15   etab = 1.847461727e-03 letab = -4.695404683e-09 wetab = -1.289832692e-09 petab = 2.579929800e-15   dsub = -1.342546866e+00 ldsub = 3.489937573e-06 wdsub = 8.547636876e-07 pdsub = -1.709702602e-12   voffl = 0.0   minv = 0.0   pclm = 4.200423067e-01 lpclm = -3.710626434e-07 wpclm = -8.844691978e-08 ppclm = 1.769119712e-13   pdiblc1 = 0.39   pdiblc2 = -7.346421110e-03 lpdiblc2 = 3.819275658e-08 wpdiblc2 = 8.768161887e-09 ppdiblc2 = -1.753812125e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.099783860e-04 lalpha0 = -5.711455483e-10 walpha0 = -1.130178786e-10 palpha0 = 2.260589259e-16   alpha1 = 0.0   beta0 = 2.728820443e+01 lbeta0 = -1.219518873e-05 wbeta0 = -3.083247051e-06 pbeta0 = 6.167126167e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.970852433e-01 lkt1 = -1.428841575e-07 wkt1 = -3.823771347e-08 pkt1 = 7.648326566e-14   kt2 = -9.696352154e-02 lkt2 = 1.197613174e-07 wkt2 = 2.470282018e-08 pkt2 = -4.941070444e-14   at = 5.245008787e+04 lat = -6.556847749e-03 wat = -1.773584866e-02 pat = 3.547533316e-8   ute = -9.627673910e-01 lute = -3.138973893e-07 wute = -9.976244042e-08 pute = 1.995453321e-13   ua1 = 2.662823072e-09 lua1 = -1.233172532e-15 wua1 = -3.072136522e-16 pua1 = 6.144902831e-22   ub1 = -2.923331619e-18 lub1 = 2.058274190e-24 wub1 = 4.671068786e-25 pub1 = -9.343095141e-31   uc1 = 4.734979477e-10 luc1 = -9.654750464e-16 wuc1 = -2.399409687e-16 puc1 = 4.799311253e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.76 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.837853312e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.257592057e-07 wvth0 = -1.277817468e-07 pvth0 = 6.391706865e-14   k1 = 2.184569275e-01 lk1 = 1.272686950e-07 wk1 = 1.214095234e-07 pk1 = -6.072965065e-14   k2 = 7.870250226e-02 lk2 = -5.943954735e-08 wk2 = -5.595224302e-08 pk2 = 2.798759172e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -9.316165088e+04 lvsat = 1.392123791e-01 wvsat = 4.135358147e-02 pvsat = -2.068526822e-8   ua = -4.440826499e-09 lua = 1.295309609e-15 wua = 1.778616719e-15 pua = -8.896729759e-22   ub = 5.786275366e-18 lub = -1.681606859e-24 wub = -1.888762106e-24 pub = 9.447682494e-31   uc = 2.270332016e-10 luc = -8.517152133e-17 wuc = -1.057317875e-16 puc = 5.288756879e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.124286274e-02 lu0 = -1.036948112e-08 wu0 = -7.663395355e-09 pu0 = 3.833268674e-15   a0 = 8.350647881e-01 la0 = 7.155693225e-08 wa0 = 5.918618603e-07 pa0 = -2.960522618e-13   keta = -4.897958542e-02 lketa = 2.449983353e-08 wketa = -9.560794975e-08 pketa = 4.782357451e-14   a1 = 0.0   a2 = 0.38689047   ags = 2.186689803e+00 lags = -9.805017425e-07 wags = 5.004521326e-07 pags = -2.503286590e-13   b0 = -1.142599305e-06 lb0 = 5.715338853e-13 wb0 = 6.203857186e-13 pb0 = -3.103200384e-19   b1 = -4.352831170e-07 lb1 = 2.177307915e-13 wb1 = 2.363413212e-13 pb1 = -1.182191106e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {4.361611021e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.325641124e-08 wvoff = -8.203304216e-08 pvoff = 4.103333785e-14   nfactor = {5.854636185e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.863640822e-06 wnfactor = -2.056261986e-06 pnfactor = 1.028552527e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.533920631e-05 lcit = 2.517992269e-11 wcit = 2.733217546e-11 pcit = -1.367169083e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.874243211e-03 leta0 = 4.181294075e-10 weta0 = -2.018929405e-09 peta0 = 1.009878583e-15   etab = -5.570077203e-03 letab = 2.723654842e-09 wetab = 2.579665384e-09 petab = -1.290361523e-15   dsub = 3.293820971e+00 ldsub = -1.147380719e-06 wdsub = -1.709527375e-06 pdsub = 8.551141407e-13   voffl = 0.0   minv = 0.0   pclm = -2.268516445e-01 lpclm = 2.759639211e-07 wpclm = 1.768938396e-07 ppclm = -8.848318302e-14   pdiblc1 = 0.39   pdiblc2 = 5.434104720e-02 lpdiblc2 = -2.350735767e-08 wpdiblc2 = -1.753632377e-08 ppdiblc2 = 8.771756834e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.630621172e-04 lalpha0 = 3.020739282e-10 walpha0 = 2.260357572e-10 palpha0 = -1.130642159e-16   alpha1 = 0.0   beta0 = 5.902823932e+00 lbeta0 = 9.194575765e-06 wbeta0 = 6.166494102e-06 pbeta0 = -3.084511182e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.092286278e-01 lkt1 = 6.930271635e-08 wkt1 = 7.647542693e-08 pkt1 = -3.825339093e-14   kt2 = 8.136751336e-02 lkt2 = -5.860627540e-08 wkt2 = -4.940564036e-08 pkt2 = 2.471294834e-14   at = 1.037861242e+04 lat = 3.552325235e-02 wat = 3.547169731e-02 pat = -1.774312035e-8   ute = -1.424061323e+00 lute = 1.474911081e-07 wute = 1.995248808e-07 pute = -9.980334302e-14   ua1 = 1.398893869e-09 lua1 = 3.101577669e-17 wua1 = 6.144273043e-16 pua1 = -3.073396098e-22   ub1 = -4.386836633e-19 lub1 = -4.268831187e-25 wub1 = -9.342137572e-25 pub1 = 4.672983924e-31   uc1 = -9.720492638e-10 luc1 = 4.803685023e-16 wuc1 = 4.798819374e-16 puc1 = -2.400393445e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.77 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.024524205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.505557715e-8   k1 = 3.451653516e-01 lk1 = 6.388850775e-8   k2 = -3.742368333e-03 lk2 = -1.820021086e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.199394048e+05 lvsat = -1.740233441e-2   ua = -1.479233181e-09 lua = -1.860941771e-16   ub = 2.549242254e-18 lub = -6.242671146e-26   uc = 7.170427229e-11 luc = -7.475214225e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.845240547e-02 lu0 = -3.971630436e-9   a0 = 4.411000044e-01 la0 = 2.686200869e-7   keta = 2.712863325e-02 lketa = -1.356987800e-8   a1 = 0.0   a2 = 0.38689047   ags = 4.531657218e-01 lags = -1.133843294e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.340416673e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.608897350e-9   nfactor = {1.667665112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.307030435e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.100000000e-09 lcit = 2.503075840e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.551186649e-03 leta0 = 7.951891478e-11   etab = 8.363960144e-03 letab = -4.246220309e-09 wetab = -1.240770919e-24 petab = -6.656013888e-31   dsub = 1.651174065e+00 ldsub = -3.257205233e-07 wdsub = -8.470329473e-22   voffl = 0.0   minv = 0.0   pclm = 9.072817740e-02 lpclm = 1.171089063e-7   pdiblc1 = 0.39   pdiblc2 = 2.372125092e-03 lpdiblc2 = 2.487757016e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.135033778e-03 lalpha0 = 6.381975126e-10 walpha0 = -2.067951531e-25   alpha1 = 0.0   beta0 = 1.863226702e+01 lbeta0 = 2.827244687e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.701295490e-01 lkt1 = -2.753383425e-10   kt2 = -4.711727502e-02 lkt2 = 5.662458166e-9   at = 1.096751699e+05 lat = -1.414538219e-02 wat = 5.551115123e-17   ute = -1.238389462e+00 lute = 5.461711484e-8   ua1 = 1.783864614e-09 lua1 = -1.615485147e-16   ub1 = -1.725425035e-18 lub1 = 2.167513493e-25   uc1 = -3.065312391e-11 luc1 = 9.477446116e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.78 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.335571740e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.435061966e-07 wvth0 = -4.136582039e-07 pvth0 = 1.034993509e-13   k1 = -2.398501938e-01 lk1 = 2.102623223e-07 wk1 = 2.748510414e-07 pk1 = -6.876910481e-14   k2 = 2.673398422e-01 lk2 = -8.602633534e-08 wk2 = -1.207576728e-07 pk2 = 3.021417352e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.155136181e+05 lvsat = 8.725519538e-03 wvsat = -1.596063585e-02 pvsat = 3.993430893e-9   ua = 3.944219775e-09 lua = -1.543069224e-15 wua = -3.286438995e-15 pua = 8.222834688e-22   ub = 7.868452908e-19 lub = 3.785338207e-25 wub = 7.000083881e-25 pub = -1.751455987e-31   uc = -2.446060692e-10 luc = 7.166721476e-17 wuc = 1.708583465e-16 puc = -4.274961258e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 9.886517055e-02 lu0 = -2.158925632e-08 wu0 = -4.941001462e-08 pu0 = 1.236263271e-14   a0 = 5.414078764e+00 la0 = -9.756440637e-7   keta = 1.501127292e+00 lketa = -3.823717123e-07 wketa = -7.238369956e-07 pketa = 1.811076355e-13   a1 = 0.0   a2 = 0.38689047   ags = -2.754147271e+00 lags = 6.891014179e-07 wags = -3.447069626e-08 pags = 8.624740557e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-6.168145325e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.264010821e-07 wvoff = 2.412542969e-07 pvoff = -6.036303135e-14   nfactor = {-6.420686258e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.254448998e-06 wnfactor = 3.858630745e-06 pnfactor = -9.654487055e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 8.765405302e-05 lcit = -1.942943233e-11 wcit = -3.517417985e-11 pcit = 8.800755670e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.030576012e-01 leta0 = 5.152386569e-08 weta0 = 1.187045559e-08 peta0 = -2.970047341e-15   etab = -1.272308973e-01 letab = 2.968029100e-08 wetab = 8.031254359e-08 petab = -2.009459997e-14   dsub = 1.067206705e-01 ldsub = 6.070943833e-08 wdsub = 1.463625763e-07 pdsub = -3.662064840e-14   voffl = 0.0   minv = 0.0   pclm = 2.247911579e+00 lpclm = -4.226291667e-07 wpclm = -4.763990919e-07 ppclm = 1.191974348e-13   pdiblc1 = -1.363150963e+01 lpdiblc1 = 3.508251818e-06 wpdiblc1 = 6.760477368e-06 ppdiblc1 = -1.691505240e-12   pdiblc2 = -1.975055184e-02 lpdiblc2 = 8.022961399e-09 wpdiblc2 = 1.449176210e-08 ppdiblc2 = -3.625911336e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.263700049e-03 lalpha0 = -7.125926846e-10 walpha0 = -2.275370561e-10 palpha0 = 5.693090913e-17   alpha1 = 0.0   beta0 = 3.731140319e+01 lbeta0 = -1.846368580e-06 wbeta0 = -1.785195150e-06 pbeta0 = 4.466647525e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 2.686257134e-01 lkt1 = -1.350745988e-07 wkt1 = -2.470634393e-07 pkt1 = 6.181650783e-14   kt2 = -1.516906248e-01 lkt2 = 3.182723316e-08 wkt2 = 6.399590283e-08 pkt2 = -1.601209487e-14   at = -5.644425546e+04 lat = 2.741852864e-02 wat = 3.029200369e-02 pat = -7.579210783e-9   ute = 1.114004543e+00 lute = -5.339636272e-07 wute = -1.252200803e-07 pute = 3.133069019e-14   ua1 = 6.707255000e-09 lua1 = -1.393405406e-15 wua1 = -1.099404166e-15 pua1 = 2.750764192e-22   ub1 = -7.516650843e-18 lub1 = 1.665745002e-24 wub1 = 1.794727353e-24 pub1 = -4.490497573e-31   uc1 = -2.147593565e-10 luc1 = 5.554174604e-17 wuc1 = 1.156920984e-16 puc1 = -2.894674149e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.79 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.439086933e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.565011696e-07 wvth0 = 9.248680578e-07 pvth0 = -1.377097741e-13   k1 = 1.972596921e+00 lk1 = -1.884317100e-07 wk1 = -6.413190966e-07 pk1 = 9.632933490e-14   k2 = -6.811572507e-01 lk2 = 8.489758329e-08 wk2 = 2.556353597e-07 pk2 = -3.761373290e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.537588509e+05 lvsat = -1.243099626e-01 wvsat = -3.392340617e-01 pvsat = 6.224891860e-8   ua = -1.473971097e-08 lua = 1.823868516e-15 wua = 6.945307256e-15 pua = -1.021528364e-21   ub = 1.903254227e-17 lub = -2.909432003e-24 wub = -8.650994329e-24 pub = 1.509951846e-30   uc = 1.490410260e-09 luc = -2.409914028e-16 wuc = -7.218182136e-16 puc = 1.181151669e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.466888615e-01 lu0 = 2.266080802e-08 wu0 = 9.357813193e-08 pu0 = -1.340454624e-14   a0 = 0.0   keta = -3.411821919e+00 lketa = 5.029663001e-07 wketa = 1.688296256e-06 pketa = -2.535708370e-13   a1 = 0.0   a2 = 0.38689047   ags = 2.023491154e-01 lags = 1.563259866e-07 wags = 8.043162460e-08 pags = -1.208123217e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {9.218619476e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.508761130e-07 wvoff = -5.629403746e-07 pvoff = 8.455686943e-14   nfactor = {1.050801041e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.961867851e-07 wnfactor = -5.907244210e-06 pnfactor = 7.944107907e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.711927904e-04 lcit = 2.721606308e-11 wcit = 8.207308633e-11 pcit = -1.232778793e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.516596662e-01 leta0 = -4.843895950e-08 weta0 = -2.769772971e-08 peta0 = 4.160337491e-15   etab = 2.354729113e-01 letab = -3.568074884e-08 wetab = -1.873959350e-07 petab = 2.814780642e-14   dsub = 1.362730394e+00 ldsub = -1.656297938e-07 wdsub = -3.415126781e-07 pdsub = 5.129691181e-14   voffl = 0.0   minv = 0.0   pclm = -8.288370269e-01 lpclm = 1.318163158e-07 wpclm = 3.915163309e-07 ppclm = -3.720526398e-14   pdiblc1 = 3.005268748e+01 lpdiblc1 = -4.363858922e-06 wpdiblc1 = -1.577444719e-05 ppdiblc1 = 2.369400840e-12   pdiblc2 = -1.010579935e-01 lpdiblc2 = 2.267496892e-08 wpdiblc2 = 5.277901273e-08 ppdiblc2 = -1.052546534e-14   pdiblcb = 0.0   drout = 7.738370796e+01 ldrout = -1.331518670e-05 wdrout = -3.346881034e-05 pdrout = 6.031246968e-12   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.777929268e-03 lalpha0 = -2.646443609e-10 walpha0 = 5.607232109e-10 palpha0 = -8.511753230e-17   alpha1 = 0.0   beta0 = 3.582160409e+01 lbeta0 = -1.577899333e-06 wbeta0 = 1.857255914e-05 pbeta0 = -3.221904359e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -8.773992193e-01 lkt1 = 7.144482423e-08 wkt1 = 3.849339196e-07 pkt1 = -5.207257622e-14   kt2 = 2.473156588e-01 lkt2 = -4.007569419e-08 wkt2 = -1.493237733e-07 pkt2 = 2.242917736e-14   at = 2.376931972e+05 lat = -2.558651103e-02 wat = -1.105095273e-01 pat = 1.779392910e-8   ute = -2.475367284e+00 lute = 1.128591229e-07 wute = 2.921801873e-07 pute = -4.388692504e-14   ua1 = -7.768521957e-09 lua1 = 1.215201980e-15 wua1 = 4.057841393e-15 pua1 = -6.542850167e-22   ub1 = 8.630035006e-18 lub1 = -1.243968521e-24 wub1 = -4.187697157e-24 pub1 = 6.290130514e-31   uc1 = 4.661629376e-10 luc1 = -6.716385596e-17 wuc1 = -2.699482297e-16 puc1 = 4.054757384e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.80 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.318901692e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.799595491e-9   k1 = 6.663443631e-01 wk1 = -6.028189310e-8   k2 = -9.450699151e-02 wk2 = 1.680421968e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.710637803e+05 wvsat = -1.225319219e-1   ua = -4.670038003e-10 wua = -2.311923692e-16   ub = 2.481904603e-18 wub = -1.490055418e-25   uc = 1.529412713e-11 wuc = 3.196294061e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.400537674e-02 wu0 = -6.971859191e-9   a0 = 2.811939279e+00 wa0 = -4.043909016e-7   keta = 3.229600000e-01 wketa = -1.462879616e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.425497094e+00 wags = 1.351328294e-6   b0 = -2.819440800e-07 wb0 = 1.277093905e-13   b1 = -1.074090431e-07 wb1 = 4.865200015e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-6.073977439e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -2.241894520e-8   nfactor = {2.147828460e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.375135196e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.785852520e-01 weta0 = -8.995117575e-8   etab = -2.439015385e-01 wetab = 7.877044086e-8   dsub = 1.305292308e+00 wdsub = -3.375876037e-7   voffl = 0.0   minv = 0.0   pclm = 8.999485538e-02 wpclm = 4.982793030e-8   pdiblc1 = 0.39   pdiblc2 = -2.159200492e-03 wpdiblc2 = 4.406530991e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -7.421626144e-05 walpha0 = 5.252125485e-11   alpha1 = 0.0   beta0 = 7.588713898e+00 wbeta0 = 4.622297857e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.628222031e-01 wkt1 = 2.351860306e-9   kt2 = -4.782162708e-02 wkt2 = 5.189846761e-9   at = -8.379257846e+03 wat = 3.017132943e-2   ute = -1.489847877e+00 wute = 1.399863263e-7   ua1 = 1.604865969e-09 wua1 = 1.624921666e-16   ub1 = -3.965055385e-19 wub1 = -4.844382113e-25   uc1 = 1.269864652e-10 wuc1 = -2.879397201e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.81 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.318901692e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.799595491e-9   k1 = 6.663443631e-01 wk1 = -6.028189310e-8   k2 = -9.450699151e-02 wk2 = 1.680421968e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.710637803e+05 wvsat = -1.225319219e-1   ua = -4.670038003e-10 wua = -2.311923692e-16   ub = 2.481904603e-18 wub = -1.490055418e-25   uc = 1.529412713e-11 wuc = 3.196294061e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.400537674e-02 wu0 = -6.971859191e-9   a0 = 2.811939279e+00 wa0 = -4.043909016e-7   keta = 3.229600000e-01 wketa = -1.462879616e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.425497094e+00 wags = 1.351328294e-6   b0 = -2.819440800e-07 wb0 = 1.277093905e-13   b1 = -1.074090431e-07 wb1 = 4.865200015e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-6.073977439e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -2.241894520e-8   nfactor = {2.147828460e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.375135196e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.785852520e-01 weta0 = -8.995117575e-8   etab = -2.439015385e-01 wetab = 7.877044086e-8   dsub = 1.305292308e+00 wdsub = -3.375876037e-7   voffl = 0.0   minv = 0.0   pclm = 8.999485538e-02 wpclm = 4.982793030e-8   pdiblc1 = 0.39   pdiblc2 = -2.159200492e-03 wpdiblc2 = 4.406530991e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -7.421626144e-05 walpha0 = 5.252125485e-11   alpha1 = 0.0   beta0 = 7.588713898e+00 wbeta0 = 4.622297857e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.628222031e-01 wkt1 = 2.351860306e-9   kt2 = -4.782162708e-02 wkt2 = 5.189846761e-9   at = -8.379257846e+03 wat = 3.017132943e-2   ute = -1.489847877e+00 wute = 1.399863263e-7   ua1 = 1.604865969e-09 wua1 = 1.624921666e-16   ub1 = -3.965055385e-19 wub1 = -4.844382113e-25   uc1 = 1.269864652e-10 wuc1 = -2.879397201e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.82 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.813607867e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.021278882e-07 wvth0 = 1.151937386e-08 pvth0 = -6.527922278e-14   k1 = 9.288441650e-01 lk1 = -1.050053020e-06 wk1 = -1.450588291e-07 pk1 = 3.391251234e-13   k2 = -1.966432426e-01 lk2 = 4.085659423e-07 wk2 = 4.979014333e-08 pk2 = -1.319504567e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.021125094e+06 lvsat = -2.200358016e+00 wvsat = -3.001797237e-01 pvsat = 7.106276248e-7   ua = -1.998263223e-11 lua = -1.788176312e-15 wua = -3.755623257e-16 pua = 5.775094216e-22   ub = 1.955051854e-18 lub = 2.107518999e-24 wub = 2.114682189e-26 pub = -6.806443360e-31   uc = -8.615984400e-11 luc = 4.058366826e-16 wuc = 3.596186858e-17 puc = -1.310690150e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.364959246e-02 lu0 = 1.423210054e-09 wu0 = -6.856955101e-09 pu0 = -4.596399190e-16   a0 = 3.136073393e+00 la0 = -1.296602904e-06 wa0 = -5.090732551e-07 pa0 = 4.187508740e-13   keta = 9.544858078e-01 lketa = -2.526232694e-06 wketa = -3.502455365e-07 pketa = 8.158721109e-13   a1 = 0.0   a2 = 0.38689047   ags = -5.343064088e+00 lags = 1.167086608e-05 wags = 2.293585730e-06 pags = -3.769222908e-12   b0 = -2.819440800e-07 wb0 = 1.277093905e-13   b1 = -1.074090431e-07 wb1 = 4.865200015e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-3.702426063e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.486691675e-08 wvoff = -3.007810752e-08 pvoff = 3.063821943e-14   nfactor = {3.822724354e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.699926929e-06 wnfactor = -6.784378975e-07 pnfactor = 2.163808401e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.556161063e-01 leta0 = -1.108180208e-06 weta0 = -1.794210605e-07 peta0 = 3.578978801e-13   etab = -4.860857444e-01 letab = 9.687864716e-07 wetab = 1.569862520e-07 petab = -3.128792789e-13   dsub = 1.855022299e+00 ldsub = -2.199032660e-06 wdsub = -5.151284017e-07 pdsub = 7.101995880e-13   voffl = 0.0   minv = 0.0   pclm = -3.033062133e-02 lpclm = 4.813265736e-07 wpclm = 8.868824626e-08 ppclm = -1.554492302e-13   pdiblc1 = 0.39   pdiblc2 = -1.672126637e-02 lpdiblc2 = 5.825124872e-08 wpdiblc2 = 9.109495786e-09 ppdiblc2 = -1.881282329e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.623978446e-04 lalpha0 = 1.152785410e-09 walpha0 = 1.455923789e-10 palpha0 = -3.723035759e-16   alpha1 = 0.0   beta0 = -4.251731170e+00 lbeta0 = 4.736420756e-05 wbeta0 = 8.446287997e-06 pbeta0 = -1.529674448e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.248742030e-01 lkt1 = -1.517997795e-07 wkt1 = -9.903825787e-09 pkt1 = 4.902525679e-14   kt2 = -4.529524507e-02 lkt2 = -1.010604593e-08 wkt2 = 4.373926429e-09 pkt2 = 3.263848592e-15   at = 2.318483622e+04 lat = -1.262628469e-01 wat = 1.997738961e-02 pat = 4.077784903e-8   ute = -1.702760898e+00 lute = 8.516957326e-07 wute = 2.087487157e-07 pute = -2.750636538e-13   ua1 = 1.316684187e-09 lua1 = 1.152786204e-15 wua1 = 2.555633548e-16 pua1 = -3.723038325e-22   ub1 = 1.095976410e-18 lub1 = -5.970233752e-24 wub1 = -9.664501813e-25 pub1 = 1.928146693e-30   uc1 = 3.800013580e-10 luc1 = -1.012111439e-15 wuc1 = -1.105076618e-16 puc1 = 3.268715103e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.83 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.478132497e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.308111605e-07 wvth0 = -4.223811359e-08 pvth0 = 4.224677241e-14   k1 = 3.280373864e-01 lk1 = 1.516837024e-07 wk1 = 4.897772808e-08 pk1 = -4.898776851e-14   k2 = 5.772295263e-02 lk2 = -1.002185932e-07 wk2 = -3.235996308e-08 pk2 = 3.236659687e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.495782885e+05 lvsat = 3.413092426e-01 wvsat = 1.102066406e-01 pvsat = -1.102292330e-7   ua = -6.450448866e-10 lua = -5.379236651e-16 wua = -1.736922200e-16 pua = 1.737278269e-22   ub = 3.997079285e-18 lub = -1.976954478e-24 wub = -6.383463571e-25 pub = 6.384772182e-31   uc = 2.083031677e-10 luc = -1.831497057e-16 wuc = -5.913790568e-17 puc = 5.915002895e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 6.630874745e-02 lu0 = -4.389974505e-08 wu0 = -1.417495580e-08 pu0 = 1.417786166e-14   a0 = 3.416067018e+00 la0 = -1.856647553e-06 wa0 = -5.994999962e-07 pa0 = 5.996228937e-13   keta = -4.870387589e-01 lketa = 3.571119518e-07 wketa = 1.153092376e-07 pketa = -1.153328760e-13   a1 = 0.0   a2 = 0.38689047   ags = -7.754179605e-01 lags = 2.534637455e-06 wags = 8.184187365e-07 pags = -8.185865124e-13   b0 = -6.774592240e-07 lb0 = 7.911113686e-13 wb0 = 2.554449614e-13 pb0 = -2.554973276e-19   b1 = -2.580839682e-07 lb1 = 3.013807386e-13 wb1 = 9.731397396e-14 pb1 = -9.733392333e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-3.873947582e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.143613475e-08 wvoff = -2.952416163e-08 pvoff = 2.953021408e-14   nfactor = {-7.760848594e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.498634254e-06 wnfactor = 8.067935261e-07 pnfactor = -8.069589188e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.101744274e-03 leta0 = -3.038218982e-09 weta0 = -9.810220928e-10 peta0 = 9.812232023e-16   etab = -3.484664834e-03 letab = 3.485379190e-09 wetab = 1.125407355e-09 petab = -1.125638063e-15   dsub = 1.251338917e+00 ldsub = -9.915421419e-07 wdsub = -3.201628168e-07 pdsub = 3.202284502e-13   voffl = 0.0   minv = 0.0   pclm = 1.763290357e-01 lpclm = 6.796489421e-08 wpclm = 2.194544342e-08 ppclm = -2.194994223e-14   pdiblc1 = 0.39   pdiblc2 = 1.331793370e-02 lpdiblc2 = -1.833309454e-09 wpdiblc2 = -5.919642686e-10 ppdiblc2 = 5.920856213e-16   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.394889233e-04 lalpha0 = -2.511320128e-10 walpha0 = -8.108897163e-11 palpha0 = 8.110559487e-17   alpha1 = 0.0   beta0 = 1.695437791e+01 lbeta0 = 4.947642146e-06 wbeta0 = 1.597563007e-06 pbeta0 = -1.597890508e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.460018991e-01 lkt1 = 9.048044378e-08 wkt1 = 2.921557493e-08 pkt1 = -2.922156412e-14   kt2 = -6.894731244e-02 lkt2 = 3.720293748e-08 wkt2 = 1.201259810e-08 pkt2 = -1.201506069e-14   at = -1.649478552e+05 lat = 2.500411031e-01 wat = 8.073672363e-02 pat = -8.075327466e-8   ute = -1.497558568e+00 lute = 4.412490055e-07 wute = 1.424765711e-07 pute = -1.425057788e-13   ua1 = 1.677992360e-09 lua1 = 4.300957921e-16 wua1 = 1.388752676e-16 pua1 = -1.389037370e-22   ub1 = -1.881167475e-18 lub1 = -1.533566844e-26 wub1 = -4.951792361e-27 pub1 = 4.952807478e-33   uc1 = -2.898685779e-10 luc1 = 3.277657561e-16 wuc1 = 1.058335327e-16 puc1 = -1.058552286e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.84 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.016815101e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.535053607e-8   k1 = 4.864927880e-01 lk1 = -6.804182572e-9   k2 = -4.482329036e-02 lk2 = 2.348671743e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.865330080e+03 lvsat = 9.354550298e-2   ua = -5.141735516e-10 lua = -6.688218288e-16   ub = 1.616454397e-18 lub = 4.041584386e-25   uc = -6.390914278e-12 luc = 3.158838857e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.432438130e-02 lu0 = -1.906772104e-9   a0 = 2.141718489e+00 la0 = -5.820377821e-7   keta = -2.600533000e-01 lketa = 1.300799609e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.291538206e+00 lags = -1.533152438e-6   b0 = 2.270265309e-07 lb0 = -1.135598059e-13   b1 = 8.648772635e-08 lb1 = -4.326159316e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.374882746e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.332907582e-9   nfactor = {1.315025654e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.070950638e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.500205000e-05 lcit = -5.003075420e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.582948165e-03 leta0 = 2.647638819e-09 weta0 = -1.033975766e-25 peta0 = 2.465190329e-32   etab = 1.250512500e-04 letab = -1.250768855e-10   dsub = -4.803034000e-01 ldsub = 7.404551622e-07 pdsub = -5.048709793e-29   voffl = 0.0   minv = 0.0   pclm = 1.636769663e-01 lpclm = 8.061955732e-8   pdiblc1 = 0.39   pdiblc2 = 1.562609715e-02 lpdiblc2 = -4.141946079e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.595712780e-05 lalpha0 = 5.246200671e-11   alpha1 = 0.0   beta0 = 1.951659579e+01 lbeta0 = 2.384899012e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.403937926e-01 lkt1 = -1.514931237e-8   kt2 = -2.770534155e-02 lkt2 = -4.047488015e-9   at = 8.868949486e+04 lat = -3.648242596e-3   ute = -9.835701520e-01 lute = -7.284477812e-8   ua1 = 2.755365311e-09 lua1 = -6.474980209e-16   ub1 = -2.501147804e-18 lub1 = 6.047717568e-25   uc1 = 8.738630976e-11 luc1 = -4.956646880e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.85 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.024524205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.505557715e-8   k1 = 3.451653516e-01 lk1 = 6.388850775e-8   k2 = -3.742368333e-03 lk2 = -1.820021086e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.199394048e+05 lvsat = -1.740233441e-2   ua = -1.479233181e-09 lua = -1.860941771e-16   ub = 2.549242254e-18 lub = -6.242671146e-26   uc = 7.170427229e-11 luc = -7.475214225e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.845240547e-02 lu0 = -3.971630436e-9   a0 = 4.411000044e-01 la0 = 2.686200869e-7   keta = 2.712863325e-02 lketa = -1.356987800e-8   a1 = 0.0   a2 = 0.38689047   ags = 4.531657218e-01 lags = -1.133843294e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.340416673e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.608897350e-9   nfactor = {1.667665112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.307030435e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -4.100000000e-09 lcit = 2.503075840e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.551186649e-03 leta0 = 7.951891478e-11   etab = 8.363960144e-03 letab = -4.246220309e-09 wetab = -4.652890946e-25 petab = 1.602373714e-31   dsub = 1.651174065e+00 ldsub = -3.257205233e-7   voffl = 0.0   minv = 0.0   pclm = 9.072817740e-02 lpclm = 1.171089063e-7   pdiblc1 = 0.39   pdiblc2 = 2.372125092e-03 lpdiblc2 = 2.487757016e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.135033778e-03 lalpha0 = 6.381975126e-10 walpha0 = 5.169878828e-26 palpha0 = -4.930380658e-32   alpha1 = 0.0   beta0 = 1.863226702e+01 lbeta0 = 2.827244687e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.701295490e-01 lkt1 = -2.753383425e-10   kt2 = -4.711727502e-02 lkt2 = 5.662458166e-9   at = 1.096751699e+05 lat = -1.414538219e-2   ute = -1.238389462e+00 lute = 5.461711484e-8   ua1 = 1.783864614e-09 lua1 = -1.615485147e-16   ub1 = -1.725425035e-18 lub1 = 2.167513493e-25 wub1 = -3.673419846e-40   uc1 = -3.065312391e-11 luc1 = 9.477446116e-18 wuc1 = 3.081487911e-33 puc1 = 7.346839693e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.86 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.223383337e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.501063207e-8   k1 = 3.669385764e-01 lk1 = 5.844073803e-8   k2 = 7.430725040e-04 lk2 = -1.932249059e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.027731501e+04 lvsat = 1.754181875e-2   ua = -3.311253104e-09 lua = 2.722863678e-16   ub = 2.332254131e-18 lub = -8.135198075e-27   uc = 1.325979808e-10 luc = -2.271112458e-17 wuc = -2.465190329e-32   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.021734142e-02 lu0 = 5.703733585e-9   a0 = 5.414078764e+00 la0 = -9.756440637e-7   keta = -9.688797590e-02 lketa = 1.745969770e-8   a1 = 0.0   a2 = 0.38689047   ags = -2.830248243e+00 lags = 7.081422616e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.419731049e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.862409944e-9   nfactor = {2.098014609e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.230274475e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.768511910e-01 leta0 = 4.496689081e-08 weta0 = 6.617444900e-24 peta0 = -7.888609052e-31   etab = 5.007514206e-02 letab = -1.468256658e-08 petab = 1.577721810e-30   dsub = 4.298453974e-01 ldsub = -2.013798397e-8   voffl = 0.0   minv = 0.0   pclm = 1.196165085e+00 lpclm = -1.594769352e-7   pdiblc1 = 1.293599357e+00 lpdiblc1 = -2.260850772e-7   pdiblc2 = 1.224291800e-02 lpdiblc2 = 1.803527681e-11   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.761366386e-03 lalpha0 = -5.869062903e-10   alpha1 = 0.0   beta0 = 3.337022704e+01 lbeta0 = -8.602666009e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.768163550e-01 lkt1 = 1.397733953e-9   kt2 = -1.040684079e-02 lkt2 = -3.522676031e-9   at = 1.043141500e+04 lat = 1.068590151e-2   ute = 8.375561143e-01 lute = -4.647948481e-7   ua1 = 4.280099919e-09 lua1 = -7.861190691e-16 pua1 = -9.403954807e-38   ub1 = -3.554430441e-18 lub1 = 6.743776469e-25 pub1 = 8.758115402e-47   uc1 = 4.065414237e-11 luc1 = -8.363988444e-18 puc1 = 7.346839693e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.87 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = -1.025e-10   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 4.852e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {4.299402e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.299402e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.076466025e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.236310864e-08 wvth0 = 8.837163580e-08 pvth0 = -1.592501063e-14   k1 = 5.567564567e-01 lk1 = 2.423460693e-8   k2 = -1.545667184e-01 lk2 = 8.665110288e-09 wk2 = 1.711091220e-08 pk2 = -3.083471934e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.921905838e+04 lvsat = 2.313867189e-02 wvsat = 2.519028267e-02 pvsat = -4.539414888e-9   ua = -3.005463693e-11 lua = -3.190020019e-16 wua = 2.824213246e-16 pua = -5.089373480e-23   ub = -4.225726033e-18 lub = 1.173645617e-24 wub = 1.884070880e-24 pub = -3.395189930e-31   uc = -3.969284417e-10 luc = 7.271218439e-17 wuc = 1.330707247e-16 puc = -2.398000995e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 5.063444232e-02 lu0 = -5.262062104e-09 wu0 = 4.198568250e-09 pu0 = -7.566029915e-16   a0 = 0.0   keta = -5.347419705e-01 lketa = 9.636317679e-08 wketa = 3.850941222e-07 pketa = -6.939588629e-14   a1 = 0.0   a2 = 0.38689047   ags = 3.799180500e-01 lags = 1.296542448e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-3.209519010e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.580195103e-08 wvoff = 4.586197739e-12 pvoff = -8.264557636e-19   nfactor = {-5.325065798e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.460703652e-06 wnfactor = 1.264505990e-06 pnfactor = -2.278703019e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.905113756e-01 leta0 = -3.925418051e-8   etab = -1.782411805e-01 letab = 2.646117632e-8   dsub = 6.087726974e-01 ldsub = -5.238157806e-8   voffl = 0.0   minv = 0.0   pclm = 3.551375667e-02 lpclm = 4.967823743e-8   pdiblc1 = -4.772566833e+00 lpdiblc1 = 8.670684012e-07 wpdiblc1 = -5.293955920e-23 ppdiblc1 = 8.204153414e-29   pdiblc2 = 1.546225717e-02 lpdiblc2 = -5.621057377e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.558925945e-03 lalpha0 = -7.306305106e-10 walpha0 = -6.989570438e-10 palpha0 = 1.259555541e-16   alpha1 = 0.0   beta0 = 1.685501616e+02 lbeta0 = -2.522036670e-05 wbeta0 = -4.154816825e-05 pbeta0 = 7.487187659e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.758042833e-02 lkt1 = -4.351582621e-8   kt2 = -8.234650400e-02 lkt2 = 9.441210978e-9   at = -1.359875667e+05 lat = 3.707133411e-02 wat = 5.875291158e-02 pat = -1.058756843e-8   ute = -1.830320950e+00 lute = 1.596993829e-8   ua1 = 2.546893904e-09 lua1 = -4.737866792e-16 wua1 = -6.146293752e-16 pua1 = 1.107592866e-22   ub1 = -6.151459300e-19 lub1 = 1.447038816e-25   uc1 = -1.298018931e-10 luc1 = 2.235304143e-17 wuc1 = -6.162975822e-33 puc1 = -7.346839693e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.49362848e-10   cgso = 2.49362848e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.408e-11   cgdl = 2.408e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.241e-9   dwc = 4.852e-8   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0013575861   mjs = 0.42197   pbs = 0.7477   cjsws = 3.62566016e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 2.01501188e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__nfet_01v8_lvt





















