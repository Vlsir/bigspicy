** Translated using xdm 2.6.0 on Nov_14_2022_16_05_35_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TOXE_MULT=1.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RSHP_MULT=1.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__OVERLAP_MULT=9.8210e-1 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AJUNCTION_MULT=1.0050e+0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PJUNCTION_MULT=1.0090e+0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__LINT_DIFF=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__WINT_DIFF=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__DLC_DIFF=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__DWC_DIFF=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_0=0.0025904 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_0=0.0013216 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_0=-5983.8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_0=0.0011957 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_0=-0.063147 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_0=1.3229e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_0=3.1718e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_0=0.019432 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_1=0.018981 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_1=0.0025296 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_1=0.0013991 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_1=-9020.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_1=0.0072841 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_1=1.4079e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_1=-0.074743 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_1=3.1631e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_2=0.016493 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_2=0.0011738 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_2=0.00094592 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_2=0.011633 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_2=-1.6818e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_2=-840.04 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_2=-0.18372 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_2=2.8322e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_3=0.020198 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_3=0.0025033 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_3=0.0015269 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_3=0.0030122 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_3=1.4317e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_3=-14143.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_3=-0.088815 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_3=2.9649e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_4=0.021723 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_4=0.0027232 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_4=0.0010803 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_4=-6.9665e-6 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_4=1.108e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_4=-2261.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_4=-0.067845 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_4=2.8628e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_5=0.022334 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_5=0.0026099 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_5=0.0013654 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_5=0.0011422 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_5=1.3711e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_5=-2378.6 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_5=-0.060725 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_5=3.6247e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_6=3.713e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_6=0.022964 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_6=0.0028181 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_6=0.0011851 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_6=0.0037406 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_6=1.6366e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_6=-232.34 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_6=-0.067505 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_7=4.2442e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_7=0.02253 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_7=0.0024309 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_7=0.0013925 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_7=0.0023129 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_7=1.816e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_7=-1157.8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_7=-0.053499 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_7=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
*




* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
.INCLUDE sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice























