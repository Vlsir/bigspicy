** Translated using xdm 2.6.0 on Nov_14_2022_16_05_06_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
.PARAM SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__TOX_SLOPE=2.0e-3
.PARAM SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_SLOPE=0.0255
.PARAM SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__TOX_SLOPE1=2.0e-3
.PARAM SKY130_FD_BS_FLASH__SPECIAL_SONOSFET_STAR__VTH0_SLOPE1=0.028
