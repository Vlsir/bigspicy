** Translated using xdm 2.6.0 on Nov_14_2022_16_05_27_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__rf_pfet_01v8_mvt_aF02W1p68L0p15 d g s b
* .param  mult = 1.0  rg_sub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult)}   rg_dist_tnom = {(250.129*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_mvt_aF02W1p68L0p15 1 2 3 b sky130_fd_pr__pfet_01v8_mvt l = 0.15 w = {(2)*(1.68)} ad = {(2)*(0.2352)} as = {(2)*(0.445)} pd = {(2)*(1.96)} ps = {(2)*(3.89)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(0.56f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(0.34f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.119f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_sub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(154*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(76*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_mvt_aF02W1p68L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15 d g s b
* .param  mult = 1.0  rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult_2)}   rg_dist_tnom = {(257.3*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult_2)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15 1 2 3 b sky130_fd_pr__pfet_01v8_mvt l = 0.15 w = {(2)*(0.84)} ad = {(2)*(0.1176)} as = {(2)*(0.223)} pd = {(2)*(1.12)} ps = {(2)*(2.21)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(0.17f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(0.300f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.100f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(306*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(152.5*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15
.SUBCKT sky130_fd_pr__rf_pfet_01v8_mvt_aF04W1p68L0p15 d g s b
* .param  mult = 1.0  rg_stub_tnom = {(88.5*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult)}   rg_dist_tnom = {(100.061*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult)}   tref = 30.0; HSpice Parser Retained (as a comment). Continuing.


* xsky130_fd_pr__rf_pfet_01v8_mvt_aF04W1p68L0p15 1 2 3 b sky130_fd_pr__pfet_01v8_mvt l = 0.15 w = {(4)*(1.68)} ad = {(4)*(0.2352)} as = {(4)*(0.34)} pd = {(4)*(1.96)} ps = {(4)*(2.925)} nrd = {(0)/(4)} nrs = {(0)/(4)} nf = 4 sa = 0.265 sb = 0.265 sd = 0.28 m = 1 mult = {1*mult}; HSpice Parser Retained (as a comment). Continuing.



* cpar_ds 1  3 c = {(0.82f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gd 2  1 c = {(0.984f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* cpar_gs 2  3 c = {(0.354f*sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}; HSpice Parser Retained (as a comment). Continuing.
* rd 1  d r = {(78*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rd_mult)}; HSpice Parser Retained (as a comment). Continuing.
* rs 3  s r = {(50.6*sky130_fd_pr__rf_pfet_01v8_mvt__aw_rs_mult)}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_pfet_01v8_mvt_aF04W1p68L0p15
