** Translated using xdm 2.6.0 on Nov_14_2022_16_05_26_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PNP_05V5_W3P40L3P40__BF_SLOPE=0.0
.PARAM SKY130_FD_PR__PNP_05V5_W3P40L3P40__IS_SLOPE=0.0
.PARAM SKY130_FD_PR__PNP_05V5_W3P40L3P40__XTI_SLOPE=0.0
*  statistics {
*   mismatch {
*     vary  sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_slope dist=gauss std=0.05537
*     vary  sky130_fd_pr__pnp_05v5_W3p40L3p40__is_slope dist=gauss std=0.01662
*     vary  sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_slope dist=gauss std=0.06
*   }
* }
.SUBCKT sky130_fd_pr__pnp_05v5_W3p40L3p40 Collector Base Emitter
* .param  mult = 1.0  sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_mm = {(16.603*dkbfpp5x*MC_MM_SWITCH*AGAUSS(0,0.05537,1)*0.45/sqrt(mult))}   sky130_fd_pr__pnp_05v5_W3p40L3p40__is_mm = {(7.1190e-018*1.00*dkispp5x*MC_MM_SWITCH*AGAUSS(0,0.01662,1)*0.13/sqrt(mult))}   sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_mm = {(5*MC_MM_SWITCH*AGAUSS(0,0.06,1)/sqrt(mult))}; HSpice Parser Retained (as a comment). Continuing.

Qsky130_fd_pr__pnp_05v5_W3p40L3p40 Collector Base Emitter Collector 
+ sky130_fd_pr__pnp_05v5_W3p40L3p40__model


* General Parameters

* Capacitance Parameters

* Noise Parameters





* DC Parameters

* Temperature Parameters






.ENDS sky130_fd_pr__pnp_05v5_W3p40L3p40


