** Translated using xdm 2.6.0 on Nov_14_2022_16_05_30_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_01V8_LVT__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_01V8_LVT__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__nfet_01v8_lvt d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__nfet_01v8_lvt d g s b sky130_fd_pr__nfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__nfet_01v8_lvt__model.0 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4171292+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.47213   k2 = -0.0343994   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 161140.0   ua = -1.3007075e-9   ub = 2.6647e-18   uc = 7.0152e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03156513   a0 = 1.9572694   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.54233   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11559919+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.0228979+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0047977   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.4345657e-5   alpha1 = 0.0   beta0 = 17.822982   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25364   kt2 = -0.034423   at = 333080.0   ute = -1.0777   ua1 = 2.6823e-9   ub1 = -2.4433e-18   uc1 = -1.9223e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.1 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.084871504e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = 6.862910821e-08 wvth0 = 6.060107626e-08 pvth0 = -4.812513269e-13   k1 = 5.482319152e-01 lk1 = -6.043481389e-07 wk1 = -5.336532648e-07 pk1 = 4.237900672e-12   k2 = -6.024068266e-02 lk2 = 2.052133780e-07 wk2 = 1.812081185e-07 pk2 = -1.439028031e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.445248009e+04 lvsat = 6.884116019e-01 wvsat = 6.078832302e-01 pvsat = -4.827383096e-6   ua = -1.338845452e-09 lua = 3.028649213e-16 wua = 2.674366705e-16 pua = -2.123794831e-21   ub = 2.669436502e-18 lub = -3.761398191e-26 wub = -3.321400855e-26 pub = 2.637624061e-31   uc = 6.984576979e-11 luc = 2.431865945e-18 wuc = 2.147393394e-18 puc = -1.705309516e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.118944170e-02 lu0 = 2.983453532e-09 wu0 = 2.634457881e-09 pu0 = -2.092102037e-14   a0 = 1.994712559e+00 la0 = -2.973473625e-07 wa0 = -2.625645395e-07 pa0 = 2.085103778e-12   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.238957892e-01 lags = 1.463915981e-07 wags = 1.292671380e-07 pags = -1.026549123e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.120979721e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.780422177e-08 wvoff = -2.455176540e-08 pvoff = 1.949729345e-13   nfactor = {1.076729949e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.274964522e-07 wnfactor = -3.774891701e-07 pnfactor = 2.997754747e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 3.393972619e-01 lpclm = -1.106995476e-06 wpclm = -9.775023893e-07 ppclm = 7.762639724e-12   pdiblc1 = 0.39   pdiblc2 = 2.901721765e-03 lpdiblc2 = 1.505653195e-08 wpdiblc2 = 1.329526297e-08 ppdiblc2 = -1.055816719e-13   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.379155021e-04 lalpha0 = -4.254142112e-10 walpha0 = -3.756505035e-10 palpha0 = 2.983153344e-15   alpha1 = 0.0   beta0 = 1.812139857e+01 lbeta0 = -2.369815497e-06 wbeta0 = -2.092601425e-06 pbeta0 = 1.661797570e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.532267482e-01 lkt1 = -3.281756811e-09 wkt1 = -2.897866517e-09 pkt1 = 2.301282737e-14   kt2 = -3.414008143e-02 lkt2 = -2.246741202e-09 wkt2 = -1.983924000e-09 pkt2 = 1.575493566e-14   at = 6.138634307e+05 lat = -2.229785458e+00 wat = -1.968951690e+00 pat = 1.563603606e-5   ute = -9.513932848e-01 lute = -1.003039518e-06 wute = -8.857068946e-07 pute = 7.033664162e-12   ua1 = 2.424812317e-09 lua1 = 2.044786936e-15 wua1 = 1.805593753e-15 pua1 = -1.433876167e-20   ub1 = -1.564027246e-18 lub1 = -6.982568723e-24 wub1 = -6.165768298e-24 pub1 = 4.896421578e-29   uc1 = -1.100564617e-11 luc1 = -6.525647198e-17 wuc1 = -5.762296114e-17 puc1 = 4.576012213e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.2 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.217756303e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.625522268e-08 wvth0 = -1.212021525e-07 pvth0 = 2.352897387e-13   k1 = 3.604411007e-01 lk1 = 1.357917983e-07 wk1 = 1.067306530e-06 pk1 = -2.071962166e-12   k2 = 2.917157061e-03 lk2 = -4.371061570e-08 wk2 = -3.624162369e-07 pk2 = 7.035586408e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.467697417e+05 lvsat = -7.790024212e-01 wvsat = -1.215766460e+00 pvsat = 2.360167430e-6   ua = -1.298795460e-09 lua = 1.450158867e-16 wua = -5.348733409e-16 pua = 1.038349617e-21   ub = 2.615527411e-18 lub = 1.748579163e-25 wub = 6.642801709e-26 pub = -1.289567096e-31   uc = 6.805343496e-11 luc = 9.495995203e-18 wuc = -4.294786787e-18 puc = 8.337469590e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.039308695e-02 lu0 = 6.122126481e-09 wu0 = -5.268915763e-09 pu0 = 1.022854617e-14   a0 = 1.854135516e+00 la0 = 2.567089394e-07 wa0 = 5.251290790e-07 pa0 = -1.019433081e-12   keta = 1.791140445e-01 lketa = -7.059421836e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.621097996e-01 lags = 3.638405425e-06 wags = -2.585342759e-07 pags = 5.018925898e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.223129836e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.245620318e-08 wvoff = 4.910353079e-08 pvoff = -9.532468432e-14   nfactor = {6.410342037e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.289711190e-06 wnfactor = 7.549783402e-07 pnfactor = -1.465639452e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 8.288957528e-01 ldsub = -1.059798831e-6   voffl = 0.0   minv = 0.0   pclm = -1.080110888e-01 lpclm = 6.563750566e-07 wpclm = 1.955004779e-06 ppclm = -3.795250777e-12   pdiblc1 = 0.39   pdiblc2 = 4.810139499e-03 lpdiblc2 = 7.534885140e-09 wpdiblc2 = -2.659052595e-08 ppdiblc2 = 5.162018802e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.301191916e-05 lalpha0 = 3.665010344e-10 walpha0 = 7.513010071e-10 palpha0 = -1.458500645e-15   alpha1 = 0.0   beta0 = 1.385447670e+01 lbeta0 = 1.444740367e-05 wbeta0 = 4.185202850e-06 pbeta0 = -8.124734294e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.544762102e-01 lkt1 = 1.642747810e-09 wkt1 = 5.795733035e-09 pkt1 = -1.125125654e-14   kt2 = -3.961689633e-02 lkt2 = 1.933902935e-08 wkt2 = 3.967848001e-09 pkt2 = -7.702783324e-15   at = 4.494718496e+04 lat = 1.248414124e-02 wat = 3.937903380e+00 pat = -7.644651832e-6   ute = -1.241498955e+00 lute = 1.403539622e-07 wute = 1.771413789e-06 pute = -3.438845589e-12   ua1 = 2.644198996e-09 lua1 = 1.180118219e-15 wua1 = -3.611187506e-15 pua1 = 7.010398306e-21   ub1 = -2.917190233e-18 lub1 = -1.649347440e-24 wub1 = 1.233153660e-23 pub1 = -2.393921199e-29   uc1 = -2.058836641e-11 luc1 = -2.748809669e-17 wuc1 = 1.152459223e-16 puc1 = -2.237269089e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.3 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.264148958e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.249016395e-9   k1 = 4.290627670e-01 lk1 = 2.576557423e-9   k2 = -1.531900303e-02 lk2 = -8.308758118e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.011825850e+04 lvsat = 4.925610307e-2   ua = -9.587073477e-10 lua = -5.151971658e-16   ub = 2.622869143e-18 lub = 1.606054127e-25   uc = 6.013673090e-11 luc = 2.486469280e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.760560307e-02 lu0 = -7.879531061e-9   a0 = 2.188489954e+00 la0 = -3.923733313e-7   keta = -1.463226330e-01 lketa = -7.417196156e-8   a1 = 0.0   a2 = 0.38689047   ags = 8.816069644e-01 lags = 1.223978071e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.170266001e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.193746774e-9   nfactor = {8.565806193e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.712709329e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.470650000e-05 lcit = -9.136728450e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.879738980e-04 leta0 = -1.707837282e-10   etab = -5.401182060e-04 letab = 7.788147331e-11   dsub = -3.965398636e-02 ldsub = 6.263167781e-7   voffl = 0.0   minv = 0.0   pclm = 2.292622430e-01 lpclm = 1.626337664e-9   pdiblc1 = 0.39   pdiblc2 = 7.074817250e-03 lpdiblc2 = 3.138466223e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.844353963e-04 lalpha0 = -1.138684391e-10   alpha1 = 0.0   beta0 = 2.120048886e+01 lbeta0 = 1.865902684e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.507872740e-01 lkt1 = -5.518583984e-9   kt2 = -4.537188610e-02 lkt2 = 3.051119099e-8   at = 3.171989080e+04 lat = 3.816228739e-2   ute = -1.318866700e+00 lute = 2.905479647e-7   ua1 = 3.273185120e-09 lua1 = -4.093254346e-17   ub1 = -3.903288500e-18 lub1 = 2.649651250e-25   uc1 = 9.639942800e-12 luc1 = -8.617031336e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.4 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.427862435e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.161333123e-9   k1 = 4.336534600e-01 lk1 = -1.744661898e-9   k2 = -2.057002668e-02 lk2 = -3.365969553e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.550509552e+04 lvsat = 4.418547339e-2   ua = -1.244279995e-09 lua = -2.463876334e-16   ub = 2.809976968e-18 lub = -1.551918298e-26   uc = 1.059038876e-10 luc = -1.821593180e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.378076078e-02 lu0 = -4.279207008e-9   a0 = 2.048208945e+00 la0 = -2.603268173e-7   keta = -4.155487592e-01 lketa = 1.792505910e-7   a1 = 0.0   a2 = 0.38689047   ags = 2.934252714e+00 lags = -7.081773726e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.149497004e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.387611347e-10   nfactor = {1.496619182e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.688026341e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 7.565262040e-04 leta0 = -3.294420138e-10   etab = -8.059310073e-04 letab = 3.280910631e-10   dsub = 2.953809615e-01 ldsub = 3.109483817e-7   voffl = 0.0   minv = 0.0   pclm = -2.145125200e-02 lpclm = 2.376229505e-7   pdiblc1 = 0.39   pdiblc2 = 1.031103140e-02 lpdiblc2 = 9.221784318e-11   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -2.148977368e-05 lalpha0 = 7.996892342e-11   alpha1 = 0.0   beta0 = 1.876746198e+01 lbeta0 = 2.476798463e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.511160980e-01 lkt1 = -5.209061953e-9   kt2 = -2.182336600e-03 lkt2 = -1.014313196e-8   at = 7.235643820e+04 lat = -8.889467766e-5   ute = -1.005433960e+00 lute = -4.486273452e-9   ua1 = 3.971613560e-09 lua1 = -6.983632340e-16   ub1 = -4.608811580e-18 lub1 = 9.290740003e-25 wub1 = 5.877471754e-39   uc1 = -1.617655314e-10 luc1 = 7.517365954e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.5 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.886299569e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.839216385e-8   k1 = 3.147669600e-01 lk1 = 5.071995055e-8   k2 = 5.158004728e-04 lk2 = -1.267114508e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.096945918e+05 lvsat = 7.032648696e-3   ua = -1.699739066e-09 lua = -4.539354531e-17   ub = 2.724306800e-18 lub = 2.228706216e-26   uc = 7.252425896e-11 luc = -3.485501679e-18 wuc = 9.860761315e-32   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.442740767e-02 lu0 = -1.515722837e-10   a0 = 1.339770520e+00 la0 = 5.230705952e-8   keta = -1.297303024e-02 lketa = 1.593921823e-9   a1 = 0.0   a2 = 0.38689047   ags = 2.346833400e+00 lags = -4.489492294e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.179930098e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.581773584e-9   nfactor = {2.070190295e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.568570188e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -4.399080946e-03 leta0 = 1.945727422e-09 weta0 = -4.394397004e-25 peta0 = 1.756448109e-31   etab = 2.078025573e-02 letab = -9.197893144e-09 wetab = -3.515517603e-24 petab = -1.035379938e-30   dsub = 1.558474961e+00 ldsub = -2.464550001e-7   voffl = 0.0   minv = 0.0   pclm = 6.217429240e-01 lpclm = -4.621863936e-8   pdiblc1 = 0.39   pdiblc2 = 7.902250800e-03 lpdiblc2 = 1.155212722e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.908797266e-03 lalpha0 = 9.128377197e-10 walpha0 = -8.271806126e-25 palpha0 = 3.451266460e-31   alpha1 = 0.0   beta0 = 1.910896638e+01 lbeta0 = 2.326092573e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.553215640e-01 lkt1 = -3.353189807e-09 wkt1 = 4.235164736e-22   kt2 = -2.786279960e-02 lkt2 = 1.189656363e-9   at = 8.511672280e+04 lat = -5.720008272e-3   ute = -5.170722000e-01 lute = -2.200003181e-7   ua1 = 3.842115324e-09 lua1 = -6.412156625e-16 wua1 = 6.310887242e-30   ub1 = -3.882137884e-18 lub1 = 6.083928982e-25   uc1 = 4.310499968e-11 luc1 = -1.523570584e-17 wuc1 = 2.465190329e-32 puc1 = 1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.6 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.832878029e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.650020979e-8   k1 = 3.743484857e-01 lk1 = 3.932200468e-8   k2 = -4.097039728e-02 lk2 = -4.734835447e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.446790886e+05 lvsat = 3.401144563e-4   ua = -1.172341397e-09 lua = -1.462847194e-16   ub = 3.085695639e-18 lub = -4.684662266e-26   uc = 7.677270943e-11 luc = -4.298230254e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.281309520e-02 lu0 = -3.668754308e-9   a0 = 4.408645143e+00 la0 = -5.347686558e-7   keta = 1.905968372e-01 lketa = -3.734899383e-08 wketa = 2.646977960e-23 pketa = 2.366582716e-29   a1 = 0.0   a2 = 0.38689047   ags = -2.086013429e+00 lags = 3.990543689e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.518953841e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.067297773e-9   nfactor = {7.242969316e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.731551023e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.184230931e-01 leta0 = 2.375852094e-08 weta0 = 3.970466940e-23 peta0 = -9.466330863e-30   etab = -4.891540181e-02 letab = 4.134886143e-9   dsub = 1.804875536e-01 ldsub = 1.715399084e-8   voffl = 0.0   minv = 0.0   pclm = 7.818336143e-01 lpclm = -7.684398841e-8   pdiblc1 = -6.670428571e-01 lpdiblc1 = 2.022122986e-7   pdiblc2 = 1.434475571e-02 lpdiblc2 = -7.723846814e-11   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 6.708847675e-03 lalpha0 = -7.357177574e-10   alpha1 = 0.0   beta0 = 3.520086395e+01 lbeta0 = -7.522874309e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.023227143e-01 lkt1 = -1.349186976e-8   kt2 = -3.211738857e-02 lkt2 = 2.003559234e-9   at = 1.237457286e+04 lat = 8.195565012e-3   ute = -1.256759429e+00 lute = -7.849815131e-8   ua1 = 1.308083120e-09 lua1 = -1.564553019e-16   ub1 = -1.708377400e-18 lub1 = 1.925525176e-25   uc1 = -1.031169707e-10 luc1 = 1.273655710e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.7 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.962270233e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = -1.167973723e-8   k1 = 9.251874667e-01 lk1 = -2.749476371e-8   k2 = -2.324406377e-01 lk2 = 1.849050472e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.707523267e+05 lvsat = -2.822569325e-3   ua = -3.134637257e-09 lua = 9.174176846e-17   ub = 3.541858277e-18 lub = -1.021791507e-25   uc = 1.464702543e-10 luc = -1.275254245e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.083583900e-02 lu0 = 2.100868693e-10   a0 = 0.0   keta = 8.148329020e-02 lketa = -2.411352057e-8   a1 = 0.0   a2 = 0.38689047   ags = 1.059850333e+00 lags = 1.746109457e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.100056323e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.986070880e-9   nfactor = {1.537025609e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.745711137e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 7.033489353e-02 leta0 = 8.621771678e-10   etab = -5.995173655e-02 letab = 5.473593547e-9   dsub = 5.103043695e-01 ldsub = -2.285278894e-8   voffl = 0.0   minv = 0.0   pclm = 1.037451667e-01 lpclm = 5.408140283e-9   pdiblc1 = 2.872891893e+00 lpdiblc1 = -2.271817866e-7   pdiblc2 = 5.069758633e-02 lpdiblc2 = -4.486836822e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.400239293e-03 lalpha0 = -9.178356065e-11   alpha1 = 0.0   beta0 = 3.062408031e+01 lbeta0 = -1.971235755e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.001897667e-01 lkt1 = -1.620596303e-9   kt2 = 1.109612000e-02 lkt2 = -3.238239356e-9   at = 6.834390000e+04 lat = 1.406485630e-3   ute = -2.583476333e+00 lute = 8.243260923e-8   ua1 = -1.755751780e-09 lua1 = 2.151878715e-16 wua1 = 2.958228395e-31   ub1 = 1.738628400e-18 lub1 = -2.255692859e-25 wub1 = -7.346839693e-40 pub1 = 4.379057701e-47   uc1 = 4.298385000e-12 luc1 = -2.929255505e-19   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.8 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.959561158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.484730768e-7   k1 = 6.585802446e-01 wk1 = -1.307454373e-6   k2 = -9.771073011e-02 wk2 = 4.439612057e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -5.124505308e+04 wvsat = 1.489318327e+0   ua = -1.394145760e-09 wua = 6.552217841e-16   ub = 2.676304464e-18 wub = -8.137456205e-26   uc = 6.940173377e-11 wuc = 5.261129403e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.064469093e-02 wu0 = 6.454440934e-9   a0 = 2.049005413e+00 wa0 = -6.432850278e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.971660498e-01 wags = 3.167054264e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.070211807e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -6.015200345e-8   nfactor = {1.154786811e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -9.248512071e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 5.415243035e-01 wpclm = -2.394887950e-6   pdiblc1 = 0.39   pdiblc2 = 1.525395615e-04 wpdiblc2 = 3.257349080e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.155921665e-04 walpha0 = -9.203464606e-10   alpha1 = 0.0   beta0 = 1.855410476e+01 wbeta0 = -5.126888683e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.526275300e-01 wkt1 = -7.099794005e-9   kt2 = -3.372984746e-02 wkt2 = -4.860628203e-9   at = 1.021001443e+06 wat = -4.823945934e+0   ute = -7.682476308e-01 wute = -2.169988321e-6   ua1 = 2.051453308e-09 wua1 = 4.423717803e-15   ub1 = -2.890753692e-19 wub1 = -1.510617709e-23   uc1 = 9.095765385e-13 wuc1 = -1.411766731e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.9 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.959561158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.484730768e-7   k1 = 6.585802446e-01 wk1 = -1.307454373e-6   k2 = -9.771073011e-02 wk2 = 4.439612057e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -5.124505308e+04 wvsat = 1.489318327e+0   ua = -1.394145760e-09 wua = 6.552217841e-16   ub = 2.676304464e-18 wub = -8.137456205e-26   uc = 6.940173377e-11 wuc = 5.261129403e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.064469093e-02 wu0 = 6.454440934e-9   a0 = 2.049005413e+00 wa0 = -6.432850278e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 4.971660498e-01 wags = 3.167054264e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.070211807e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -6.015200345e-8   nfactor = {1.154786811e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -9.248512071e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 5.415243035e-01 wpclm = -2.394887950e-6   pdiblc1 = 0.39   pdiblc2 = 1.525395615e-04 wpdiblc2 = 3.257349080e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.155921665e-04 walpha0 = -9.203464606e-10   alpha1 = 0.0   beta0 = 1.855410476e+01 wbeta0 = -5.126888683e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.526275300e-01 wkt1 = -7.099794004e-9   kt2 = -3.372984746e-02 wkt2 = -4.860628203e-9   at = 1.021001443e+06 wat = -4.823945934e+0   ute = -7.682476308e-01 wute = -2.169988321e-6   ua1 = 2.051453308e-09 wua1 = 4.423717803e-15   ub1 = -2.890753692e-19 wub1 = -1.510617709e-23   uc1 = 9.095765385e-13 wuc1 = -1.411766731e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.10 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.574087676e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.519266637e-07 wvth0 = 3.301608170e-07 pvth0 = -7.160858906e-13   k1 = 1.043613452e+00 lk1 = -1.517531379e-06 wk1 = -3.723337105e-06 pk1 = 9.521718614e-12   k2 = -2.311112020e-01 lk2 = 5.257712800e-07 wk2 = 1.278672527e-06 pk2 = -3.289847731e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.372672715e+05 lvsat = 3.390393696e-01 wvsat = 2.879705489e+00 pvsat = -5.479932922e-6   ua = -1.626428165e-09 lua = 9.154946406e-16 wua = 1.762601855e-15 pua = -4.364517073e-21   ub = 2.584216531e-18 lub = 3.629461709e-25 wub = 2.859908710e-25 pub = -1.447897381e-30   uc = 1.248621858e-10 luc = -2.185862796e-16 wuc = -4.026576307e-16 puc = 1.607730209e-21   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.498401150e-02 lu0 = 2.231043582e-08 wu0 = 3.266141448e-08 pu0 = -1.032895448e-13   a0 = 1.958838801e+00 la0 = 3.553736647e-07 wa0 = -2.090870050e-07 pa0 = -1.711304667e-12   keta = 9.981335590e-02 lketa = -3.933943796e-07 wketa = 5.560841837e-07 pketa = -2.191694593e-12   a1 = 0.0   a2 = 0.38689047   ags = -7.219856279e-01 lags = 4.805042507e-06 wags = 2.265040988e-06 pags = -7.678974950e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.695103593e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.910246164e-08 wvoff = -1.988668232e-07 pvoff = 5.467167189e-13   nfactor = {1.240255398e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.368573419e-07 wnfactor = -3.446970404e-06 pnfactor = 9.940428390e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -2.599410327e-06 lcit = 4.965805592e-11 wcit = 8.835147501e-11 pcit = -3.482196684e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 1.177604593e+00 ldsub = -2.434164981e-06 wdsub = -2.445268433e-06 pdsub = 9.637536476e-12   voffl = 0.0   minv = 0.0   pclm = 3.882287456e-01 lpclm = 6.041837823e-07 wpclm = -1.524802624e-06 ppclm = -3.429267295e-12   pdiblc1 = 0.39   pdiblc2 = -7.904225226e-03 lpdiblc2 = 3.175412706e-08 wpdiblc2 = 6.256704954e-08 ppdiblc2 = -1.182136130e-13   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.111312108e-04 lalpha0 = -3.765480355e-10 walpha0 = -1.872321570e-09 palpha0 = 3.752019500e-15   alpha1 = 0.0   beta0 = 1.594451045e+01 lbeta0 = 1.028519406e-05 wbeta0 = -1.047084532e-05 pbeta0 = 2.106213629e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.792975888e-01 lkt1 = 1.051147026e-07 wkt1 = 1.798519271e-07 pkt1 = -7.368328184e-13   kt2 = -1.801237887e-02 lkt2 = -6.194725898e-08 wkt2 = -1.475305900e-07 pkt2 = 5.623051206e-13   at = 1.979432671e+06 lat = -3.777464996e+00 wat = -9.627385916e+00 pat = 1.893179800e-5   ute = -5.408396422e-01 lute = -8.962831055e-07 wute = -3.141854546e-06 pute = 3.830416353e-12   ua1 = -6.825809899e-10 lua1 = 1.077564938e-14 wua1 = 1.971735813e-14 pua1 = -6.027682461e-20   ub1 = 5.332548929e-18 lub1 = -2.215650784e-23 wub1 = -4.551852182e-23 pub1 = 1.198641743e-28   uc1 = 2.354864351e-11 luc1 = -8.922735467e-17 wuc1 = -1.942582393e-16 puc1 = 2.092103768e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.11 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.308292513e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.395478672e-09 wvth0 = -3.095500529e-08 pvth0 = -1.505174475e-14   k1 = 1.112436494e-01 lk1 = 2.924781183e-07 wk1 = 2.228658889e-06 pk1 = -2.032891210e-12   k2 = 9.746324346e-02 lk2 = -1.120902910e-07 wk2 = -7.908685862e-07 pk2 = 7.277524323e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.146936014e+03 lvsat = 5.674676851e-02 wvsat = 8.394710323e-02 pvsat = -5.252716775e-8   ua = -8.836762589e-10 lua = -5.264096341e-16 wua = -5.261442559e-16 pua = 7.862575178e-23   ub = 2.660441391e-18 lub = 2.149708502e-25 wub = -2.634697510e-25 pub = -3.812294759e-31   uc = -8.302818911e-11 luc = 1.849913052e-16 wuc = 1.003922527e-15 puc = -1.122863851e-21   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.167675071e-02 lu0 = -1.009517881e-08 wu0 = -2.854831217e-08 pu0 = 1.553689751e-14   a0 = 2.476009631e+00 la0 = -6.486100675e-07 wa0 = -2.016188609e-06 pa0 = 1.796821677e-12   keta = 1.491496647e-01 lketa = -4.891709559e-07 wketa = -2.071955167e-06 pketa = 2.910118198e-12   a1 = 0.0   a2 = 0.38689047   ags = 9.485518252e-01 lags = 1.562028149e-06 wags = -4.694407944e-07 pags = -2.370525465e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.420307204e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.782372982e-08 wvoff = 1.753376432e-07 pvoff = -1.797264116e-13   nfactor = {5.964651091e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.955058691e-06 wnfactor = 5.588380895e-06 pnfactor = -7.599899087e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 3.990532065e-05 lcit = -3.285637833e-11 wcit = -1.767029500e-10 pcit = 1.663304868e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 7.493794381e-04 leta0 = -4.841203031e-10 weta0 = -1.131832139e-09 peta0 = 2.197225731e-15   etab = -5.864016417e-04 letab = 1.677315071e-10 wetab = 3.245556504e-10 petab = -6.300598842e-16   dsub = 1.775509467e-01 ldsub = -4.927608381e-07 wdsub = -1.523117012e-06 pdsub = 7.847363922e-12   voffl = 0.0   minv = 0.0   pclm = 1.244033697e+00 lpclm = -1.057190369e-06 wpclm = -7.115932605e-06 ppclm = 7.424793336e-12   pdiblc1 = 0.39   pdiblc2 = 1.056554883e-02 lpdiblc2 = -4.101245314e-09 wpdiblc2 = -2.447823158e-08 ppdiblc2 = 5.076739120e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.587633762e-04 lalpha0 = -8.075635811e-11 walpha0 = 1.800211900e-10 palpha0 = -2.321935008e-16   alpha1 = 0.0   beta0 = 2.069638527e+01 lbeta0 = 1.060379475e-06 wbeta0 = 3.534950813e-06 pbeta0 = -6.127315741e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.144885111e-01 lkt1 = -2.069915991e-08 wkt1 = -2.545396301e-07 pkt1 = 1.064515116e-13   kt2 = -1.401206010e-01 lkt2 = 1.751014327e-07 wkt2 = 6.644111512e-07 pkt2 = -1.013917382e-12   at = 8.358519771e+02 lat = 6.358500813e-02 wat = 2.165696896e-01 pat = -1.782730158e-7   ute = -1.392657383e+00 lute = 7.573506744e-07 wute = 5.174460944e-07 pute = -3.273383981e-12   ua1 = 3.836502556e-09 lua1 = 2.002752490e-15 wua1 = -3.950179019e-15 pua1 = -1.433103475e-20   ub1 = -4.821582097e-18 lub1 = -2.444293284e-24 wub1 = 6.439396107e-24 pub1 = 1.899826821e-29   uc1 = 1.650640087e-10 luc1 = -3.639511331e-16 wuc1 = -1.089887949e-15 puc1 = 1.947896331e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.12 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.514797635e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.004284850e-08 wvth0 = -6.096200528e-08 pvth0 = 1.319384434e-14   k1 = 4.478729521e-01 lk1 = -2.439104436e-08 wk1 = -9.971205564e-08 pk1 = 1.588043600e-13   k2 = -3.113185648e-02 lk2 = 8.956276544e-09 wk2 = 7.406324718e-08 pk2 = -8.640790242e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.254316887e+05 lvsat = -5.365336923e-02 wvsat = -7.007202460e-01 pvsat = 6.860802081e-7   ua = -6.981000185e-10 lua = -7.010925491e-16 wua = -3.830005155e-15 pua = 3.188550016e-21   ub = 2.518625548e-18 lub = 3.484621031e-25 wub = 2.043058131e-24 pub = -2.552364171e-30   uc = 1.364856405e-10 luc = -2.163706256e-17 wuc = -2.144499548e-16 puc = 2.399016632e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.878055858e-02 lu0 = -7.368993159e-09 wu0 = -3.506033215e-08 pu0 = 2.166666192e-14   a0 = 2.321730589e+00 la0 = -5.033872051e-07 wa0 = -1.918029503e-06 pa0 = 1.704424510e-12   keta = -6.678414158e-01 lketa = 2.798627482e-07 wketa = 1.769164411e-06 pketa = -7.055276607e-13   a1 = 0.0   a2 = 0.38689047   ags = 8.092530099e-01 lags = 1.693150124e-06 wags = 1.490124167e-05 pags = -1.683894887e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.109463908e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.435949632e-09 wvoff = -2.807260821e-08 pvoff = 1.174365805e-14   nfactor = {2.940861630e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.570291007e-07 wnfactor = -1.012753353e-05 pnfactor = 7.193491165e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.108021900e-04 leta0 = -1.654175009e-10 weta0 = 2.424338077e-09 peta0 = -1.150197293e-15   etab = -7.147974272e-04 letab = 2.885904599e-10 wetab = -6.390605602e-10 petab = 2.769920549e-16   dsub = -1.533864264e+00 ldsub = 1.118194300e-06 wdsub = 1.282730776e-05 pdsub = -5.660690913e-12   voffl = 0.0   minv = 0.0   pclm = -5.319062373e-01 lpclm = 6.145018906e-07 wpclm = 3.579489016e-06 ppclm = -2.642807036e-12   pdiblc1 = 0.39   pdiblc2 = 9.565343593e-04 lpdiblc2 = 4.943720006e-09 wpdiblc2 = 6.559700732e-08 ppdiblc2 = -3.402043119e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -9.543529085e-05 lalpha0 = 1.585208472e-10 walpha0 = 5.185318473e-10 palpha0 = -5.508335825e-16   alpha1 = 0.0   beta0 = 1.855749810e+01 lbeta0 = 3.073713969e-06 wbeta0 = 1.472340280e-06 pbeta0 = -4.185780446e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.191902242e-01 lkt1 = -1.627343738e-08 wkt1 = -2.238754013e-07 pkt1 = 7.758727305e-14   kt2 = 8.741138396e-02 lkt2 = -3.907442475e-08 wkt2 = -6.282625264e-07 pkt2 = 2.028763510e-13   at = 1.490308609e+04 lat = 5.034352066e-02 wat = 4.028830137e-01 pat = -3.536497477e-7   ute = -2.771945073e-01 lute = -2.926345303e-07 wute = -5.106669926e-06 pute = 2.020596429e-12   ua1 = 9.154541883e-09 lua1 = -3.003117929e-15 wua1 = -3.634450743e-14 pua1 = 1.616174658e-20   ub1 = -1.187204758e-17 lub1 = 4.192309873e-24 wub1 = 5.093235295e-23 pub1 = -2.288295207e-29   uc1 = -5.040881209e-10 luc1 = 2.659217665e-16 wuc1 = 2.400485811e-15 puc1 = -1.337592488e-21   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.13 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.838790107e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.434063627e-08 wvth0 = 3.331529767e-08 pvth0 = -2.841072945e-14   k1 = 2.916541079e-01 lk1 = 4.454833159e-08 wk1 = 1.620754083e-07 pk1 = 4.327755222e-14   k2 = 1.862885136e-02 lk2 = -1.300312383e-08 wk2 = -1.270150524e-07 pk2 = 2.327951172e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.085381786e+05 lvsat = 4.959753322e-02 wvsat = 1.530324567e+00 pvsat = -2.984798680e-7   ua = -2.071118832e-09 lua = -9.517934674e-17 wua = 2.604244904e-15 pua = 3.491154647e-22   ub = 3.330693629e-18 lub = -9.903541283e-27 wub = -4.252196683e-24 pub = 2.257317781e-31   uc = 1.281726996e-10 luc = -1.796856175e-17 wuc = -3.902263426e-16 puc = 1.015602863e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.547006903e-02 lu0 = -1.495074119e-09 wu0 = -7.311506366e-09 pu0 = 9.421105096e-15   a0 = 5.187995112e-01 la0 = 2.922462796e-07 wa0 = 5.756936054e-06 pa0 = -1.682537790e-12   keta = -1.169425109e-01 lketa = 3.675106146e-08 wketa = 7.290703875e-07 pketa = -2.465341681e-13   a1 = 0.0   a2 = 0.38689047   ags = 8.201093910e+00 lags = -1.568869265e-06 wags = -4.105212369e-05 pags = 7.853271262e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.218475152e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.374716558e-09 wvoff = 2.702914049e-08 pvoff = -1.257274366e-14   nfactor = {9.188254925e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.352954469e-07 wnfactor = 8.073772972e-06 pnfactor = -8.387453957e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -8.697354342e-03 leta0 = 3.854012342e-09 weta0 = 3.014100355e-08 peta0 = -1.338156177e-14   etab = -3.671704426e-02 letab = 1.617638199e-08 wetab = 4.031911916e-07 petab = -1.779332982e-13   dsub = 1.696224275e+00 ldsub = -3.072437725e-07 wdsub = -9.659464035e-07 pdsub = 4.262721479e-13   voffl = 0.0   minv = 0.0   pclm = 1.252717177e+00 lpclm = -1.730524222e-07 wpclm = -4.424612304e-06 ppclm = 8.894028771e-13   pdiblc1 = 0.39   pdiblc2 = 1.273255638e-02 lpdiblc2 = -2.530385136e-10 wpdiblc2 = -3.387179336e-08 ppdiblc2 = 9.875150552e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.749714036e-03 lalpha0 = 1.771154057e-09 walpha0 = 1.290915271e-08 palpha0 = -6.018814571e-15   alpha1 = 0.0   beta0 = 1.959375109e+01 lbeta0 = 2.616415523e-06 wbeta0 = -3.399480046e-06 pbeta0 = -2.035846137e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.892100871e-01 lkt1 = -2.950367185e-08 wkt1 = -4.635968147e-07 pkt1 = 1.833763328e-13   kt2 = 6.026796657e-03 lkt2 = -3.159406373e-09 wkt2 = -2.376457103e-07 pkt2 = 3.049715008e-14   at = 1.724021416e+05 lat = -1.916081252e-02 wat = -6.120759063e-01 pat = 9.425162367e-8   ute = 1.259984593e+00 lute = -9.709916674e-07 wute = -1.246134420e-05 pute = 5.266214188e-12   ua1 = 7.837947194e-09 lua1 = -2.422104692e-15 wua1 = -2.802017161e-14 pua1 = 1.248821719e-20   ub1 = -6.958546162e-18 lub1 = 2.023981698e-24 wub1 = 2.157285159e-23 pub1 = -9.926604119e-30   uc1 = 2.744129895e-10 luc1 = -7.763077353e-17 wuc1 = -1.622012583e-15 puc1 = 4.375360529e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.14 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.672041754e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.028074029e-08 wvth0 = 1.127840247e-07 pvth0 = -4.361309694e-14   k1 = 2.459613929e-01 lk1 = 5.328934797e-08 wk1 = 9.002952302e-07 pk1 = -9.794389972e-14   k2 = 2.203351484e-02 lk2 = -1.365443595e-08 wk2 = -4.418054832e-07 pk2 = 6.254736059e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.600657509e+05 lvsat = -1.786398499e-03 wvsat = -1.078966618e-01 pvsat = 1.491185312e-8   ua = -2.909809034e-09 lua = 6.526208894e-17 wua = 1.218373119e-14 pua = -1.483440261e-21   ub = 4.585981213e-18 lub = -2.500400561e-25 wub = -1.052052755e-23 pub = 1.424863473e-30   uc = -3.272731127e-12 luc = 7.176949147e-18 wuc = 5.613066451e-16 puc = -8.046797427e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.943740287e-02 lu0 = -2.254025084e-09 wu0 = 9.379503609e-08 pu0 = -9.920576475e-15   a0 = 5.592751802e+00 la0 = -6.784007935e-07 wa0 = -8.303370329e-06 pa0 = 1.007198821e-12   keta = 5.567418731e-01 lketa = -9.212476119e-08 wketa = -2.567537142e-06 pketa = 3.841068522e-13   a1 = 0.0   a2 = 0.38689047   ags = -2.139547131e+00 lags = 4.092953661e-07 wags = 3.753970568e-07 pags = -7.181345697e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.589935552e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.048075401e-08 wvoff = 4.977486004e-08 pvoff = -1.692399981e-14   nfactor = {-4.483037875e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.968272782e-07 wnfactor = 8.222686652e-06 pnfactor = -8.672325828e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 8.843055796e-07 lcit = 7.873323426e-13 wcit = 2.886068977e-11 pcit = -5.521049953e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -4.206297472e-02 leta0 = 1.023685535e-08 weta0 = -5.354638760e-07 peta0 = 9.481865170e-14   etab = 1.467078980e-01 letab = -1.891280947e-08 wetab = -1.371779046e-06 petab = 1.616185083e-13   dsub = -3.291179115e-01 ldsub = 8.020418775e-08 wdsub = 3.573531883e-06 pdsub = -4.421300483e-13   voffl = 0.0   minv = 0.0   pclm = 6.443051412e-01 lpclm = -5.666319974e-08 wpclm = 9.643977879e-07 ppclm = -1.415147534e-13   pdiblc1 = -6.670494251e-01 lpdiblc1 = 2.022135550e-07 wpdiblc1 = 4.605711790e-11 ppdiblc1 = -8.810726654e-18   pdiblc2 = -8.637193264e-03 lpdiblc2 = 3.834994594e-09 wpdiblc2 = 1.611574699e-07 ppdiblc2 = -2.743394751e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.768063066e-02 lalpha0 = -2.328470884e-09 walpha0 = -7.693798245e-08 palpha0 = 1.116894239e-14   alpha1 = 0.0   beta0 = 4.692999869e+01 lbeta0 = -2.613008642e-06 wbeta0 = -8.224879800e-05 pbeta0 = 1.304802839e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.745790938e-01 lkt1 = 5.957419113e-09 wkt1 = 1.207922023e-06 pkt1 = -1.363852208e-13   kt2 = -7.181456452e-02 lkt2 = 1.173164602e-08 wkt2 = 2.783704918e-07 pkt2 = -6.821674938e-14   at = 7.284741810e+04 lat = -1.159939214e-04 wat = -4.240567564e-01 pat = 5.828356029e-8   ute = -5.711696336e+00 lute = 3.626908943e-07 wute = 3.123957682e-05 pute = -3.093772004e-12   ua1 = -1.199915966e-08 lua1 = 1.372733848e-15 wua1 = 9.331504388e-14 pua1 = -1.072320953e-20   ub1 = 9.888346947e-18 lub1 = -1.198828954e-24 wub1 = -8.132028998e-23 pub1 = 9.756853863e-30   uc1 = -3.708165588e-10 luc1 = 4.580163906e-17 wuc1 = 1.877203206e-15 puc1 = -2.318639275e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.15 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.05e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.559560126e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.678633814e-08 wvth0 = -1.120075578e-06 pvth0 = 1.059327729e-13   k1 = 1.346013440e+00 lk1 = -8.014696530e-08 wk1 = -2.950979012e-06 pk1 = 3.692156658e-13   k2 = -3.680460443e-01 lk2 = 3.366221457e-08 wk2 = 9.509125723e-07 pk2 = -1.063893395e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.066899662e+05 lvsat = 4.688084186e-03 wvsat = 4.492276933e-01 pvsat = -5.266733115e-8   ua = -5.901832385e-09 lua = 4.281945214e-16 wua = 1.940454076e-14 pua = -2.359324462e-21   ub = 6.840962349e-18 lub = -5.235692679e-25 wub = -2.313447244e-23 pub = 2.954934989e-30   uc = 3.147042971e-10 luc = -3.139366437e-17 wuc = -1.179715990e-15 puc = 1.307180713e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.825537215e-03 lu0 = 9.739942208e-10 wu0 = 5.617103972e-08 pu0 = -5.356785716e-15   a0 = 0.0   keta = 3.804170026e-01 lketa = -7.073655440e-08 wketa = -2.096227818e-06 pketa = 3.269370313e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.190292814e+00 lags = 5.385780768e-09 wags = -9.147083322e-07 pags = 8.467632671e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-3.265205664e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.080178047e-08 wvoff = 1.518278498e-06 pvoff = -1.950534911e-13   nfactor = {-1.223849075e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.909009216e-07 wnfactor = 1.936021959e-05 pnfactor = -2.218215328e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.460328698e-05 lcit = -8.767801014e-13 wcit = -6.734160946e-11 pcit = 6.148288944e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.174671772e-01 leta0 = 3.151338511e-08 weta0 = 2.018168850e-06 peta0 = -2.149369980e-13   etab = -1.308046486e-01 letab = 1.474946243e-08 wetab = 4.968454175e-07 petab = -6.504563916e-14   dsub = 5.514728362e-01 ldsub = -2.661146994e-08 wdsub = -2.886876974e-07 pdsub = 2.635718678e-14   voffl = 0.0   minv = 0.0   pclm = 1.053733393e+00 lpclm = -1.063268467e-07 wpclm = -6.661649939e-06 ppclm = 7.835248358e-13   pdiblc1 = 6.844952824e+00 lpdiblc1 = -7.089923177e-07 wpdiblc1 = -2.785348147e-05 ppdiblc1 = 3.378624078e-12   pdiblc2 = 9.905544587e-02 lpdiblc2 = -9.228122533e-09 wpdiblc2 = -3.391022363e-07 ppdiblc2 = 3.324755485e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.340780696e-03 lalpha0 = 4.640263143e-10 walpha0 = 4.727039152e-08 palpha0 = -3.897533377e-15   alpha1 = 0.0   beta0 = 2.158819392e+01 lbeta0 = 4.609522758e-07 wbeta0 = 6.336279791e-05 pbeta0 = -4.614658196e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.946281552e-02 lkt1 = -3.711818544e-08 wkt1 = -1.968555636e-06 pkt1 = 2.489215192e-13   kt2 = 2.730312039e-01 lkt2 = -3.009814569e-08 wkt2 = -1.836780486e-06 pkt2 = 1.883510642e-13   at = -3.745173830e+04 lat = 1.326329375e-02 wat = 7.418760442e-01 pat = -8.314408842e-8   ute = -3.863433119e+00 lute = 1.384965662e-07 wute = 8.975504967e-06 pute = -3.931400883e-13   ua1 = -5.211686798e-09 lua1 = 5.494133903e-16 wua1 = 2.423422592e-14 pua1 = -2.343706317e-21   ub1 = 4.362349735e-18 lub1 = -5.285254921e-25 wub1 = -1.839845230e-23 pub1 = 2.124434952e-30   uc1 = -1.885078564e-10 luc1 = 2.368759346e-17 wuc1 = 1.352024847e-15 puc1 = -1.681597925e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.16 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.425285+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40031   k2 = -0.010012091   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 242950.0   ua = -1.2647154e-9   ub = 2.66023e-18   uc = 7.0441e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03191968   a0 = 1.921933   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.559727   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.97209474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.068446   pdiblc1 = 0.39   pdiblc2 = 0.006587   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.3789948e-5   alpha1 = 0.0   beta0 = 17.541356   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25403   kt2 = -0.03469   at = 68095.0   ute = -1.1969   ua1 = 2.9253e-9   ub1 = -3.2731e-18   uc1 = -2.6978e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.17 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.425285+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40031   k2 = -0.010012091   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 242950.0   ua = -1.2647154e-9   ub = 2.66023e-18   uc = 7.0441e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03191968   a0 = 1.921933   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.559727   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.97209474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.068446   pdiblc1 = 0.39   pdiblc2 = 0.006587   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.3789948e-5   alpha1 = 0.0   beta0 = 17.541356   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25403   kt2 = -0.03469   at = 68095.0   ute = -1.1969   ua1 = 2.9253e-9   ub1 = -3.2731e-18   uc1 = -2.6978e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.18 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.226276515e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.047340766e-8   k1 = 3.081176630e-01 lk1 = 3.633576578e-7   k2 = 2.147357124e-02 lk2 = -1.240944406e-07 pk2 = 3.231174268e-27   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.315802971e+05 lvsat = -7.434485900e-1   ua = -1.278249581e-09 lua = 5.334226609e-17   ub = 2.640710228e-18 lub = 7.693327541e-26   uc = 4.532251930e-11 luc = 9.899946798e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.143584009e-02 lu0 = 1.906958220e-9   a0 = 1.917536441e+00 la0 = 1.732815868e-8   keta = 2.096604000e-01 lketa = -8.263345345e-7   a1 = 0.0   a2 = 0.38689047   ags = -2.745568668e-01 lags = 3.288163004e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.262345353e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.889416422e-8   nfactor = {5.593521806e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.626742249e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.485325000e-05 lcit = -1.912811423e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 6.945742939e-01 ldsub = -5.303976644e-7   voffl = 0.0   minv = 0.0   pclm = 8.702424100e-02 lpclm = -7.322242125e-8   pdiblc1 = 0.39   pdiblc2 = 4.455064340e-03 lpdiblc2 = 8.402598017e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.872104563e-05 lalpha0 = 3.646135792e-10 palpha0 = 1.262177448e-29   alpha1 = 0.0   beta0 = 1.387613404e+01 lbeta0 = 1.444573932e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.437702295e-01 lkt1 = -4.043683347e-8   kt2 = -4.715508730e-02 lkt2 = 4.912864858e-8   at = 7.767046225e+04 lat = -3.773976937e-2   ute = -1.161471275e+00 lute = -1.396352338e-7   ua1 = 3.212321205e-09 lua1 = -1.131236675e-15   ub1 = -3.659030440e-18 lub1 = 1.521067643e-24   uc1 = -1.482449135e-11 luc1 = -4.790062364e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.19 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.247145012e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.422206428e-9   k1 = 5.514856100e-01 lk1 = -1.090925377e-7   k2 = -5.876234074e-02 lk2 = 3.166753534e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.472957120e+04 lvsat = 4.637072423e-2   ua = -9.876090679e-10 lua = -5.108781612e-16   ub = 2.608396441e-18 lub = 1.396640311e-25   uc = 1.152833711e-10 luc = -3.681553362e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.603741085e-02 lu0 = -7.026071084e-9   a0 = 2.077738352e+00 la0 = -2.936718122e-07 wa0 = 2.168404345e-19   keta = -2.601375570e-01 lketa = 8.568423940e-8   a1 = 0.0   a2 = 0.38689047   ags = 8.558200317e-01 lags = 1.093762331e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.073950980e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.678835512e-9   nfactor = {1.163556927e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.537995750e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.258010330e-04 leta0 = -5.008754536e-11   etab = -5.222899840e-04 letab = 4.327154594e-11   dsub = -1.233205877e-01 ldsub = 1.057381669e-06 pdsub = -5.169878828e-26   voffl = 0.0   minv = 0.0   pclm = -1.616242692e-01 lpclm = 4.094789316e-07 ppclm = -1.292469707e-26   pdiblc1 = 0.39   pdiblc2 = 5.730199320e-03 lpdiblc2 = 5.927178480e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.943241711e-04 lalpha0 = -1.266231000e-10   alpha1 = 0.0   beta0 = 2.139466785e+01 lbeta0 = -1.499903616e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.647694340e-01 lkt1 = 3.289222242e-10   kt2 = -8.875003400e-03 lkt2 = -2.518447830e-8   at = 4.361631750e+04 lat = 2.836954184e-2   ute = -1.290442780e+00 lute = 1.107371488e-7   ua1 = 3.056197160e-09 lua1 = -8.281530667e-16   ub1 = -3.549564930e-18 lub1 = 1.308562249e-24 wub1 = 3.761581923e-37   uc1 = -5.022887870e-11 luc1 = 2.082991352e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.20 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.394375291e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.436579801e-9   k1 = 4.281761600e-01 lk1 = 6.978647592e-9   k2 = -1.650164577e-02 lk2 = -8.112456835e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -1.298628828e+04 lvsat = 8.187266276e-2   ua = -1.454666663e-09 lua = -7.123684659e-17   ub = 2.922204544e-18 lub = -1.557235363e-25   uc = 9.412390042e-11 luc = -1.689812386e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.185485567e-02 lu0 = -3.089031893e-09 wu0 = -3.388131789e-21   a0 = 1.942849338e+00 la0 = -1.667007828e-7   keta = -3.183664860e-01 lketa = 1.404951303e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.752795371e+00 lags = -1.633160556e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.164917617e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.838540254e-10   nfactor = {9.403019033e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.639495289e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.896980230e-04 leta0 = -3.926236983e-10   etab = -8.410353523e-04 letab = 3.433065611e-10   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 1.751742720e-01 lpclm = 9.245046477e-8   pdiblc1 = 0.39   pdiblc2 = 1.391435184e-02 lpdiblc2 = -1.776564287e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 6.993788002e-06 lalpha0 = 4.971098959e-11   alpha1 = 0.0   beta0 = 1.884833936e+01 lbeta0 = 2.246868641e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.634138360e-01 lkt1 = -9.471021732e-10   kt2 = -3.669353300e-02 lkt2 = 1.001103613e-9   at = 9.448727400e+04 lat = -1.951528952e-2   ute = -1.285949320e+00 lute = 1.065074549e-7   ua1 = 1.975167200e-09 lua1 = 1.894204346e-16   ub1 = -1.811037780e-18 lub1 = -3.279133577e-25   uc1 = -2.990403440e-11 luc1 = 1.698137581e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.21 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.289304675e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.295901865e-07 wvth0 = 1.830189055e-06 pvth0 = -8.076624301e-13   k1 = 3.236699520e-01 lk1 = 5.309723718e-8   k2 = 2.230459153e-02 lk2 = -2.523764936e-08 wk2 = -1.456229357e-07 pk2 = 6.426340151e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.119086049e+05 lvsat = 2.675654641e-02 wvsat = 4.143457929e-01 pvsat = -1.828507984e-7   ua = -3.478681877e-09 lua = 8.219610674e-16 wua = 9.729821687e-15 pua = -4.293770311e-21   ub = 4.936978806e-18 lub = -1.044843418e-24 wub = -1.238377445e-23 pub = 5.464959664e-30   uc = 5.108866892e-11 luc = 2.093323795e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.305408916e-02 lu0 = 5.207746365e-09 wu0 = 5.554252930e-08 pu0 = -2.451091818e-14   a0 = 1.656005760e+00 la0 = -4.011671189e-8   keta = 2.707566004e-02 lketa = -1.194848878e-8   a1 = 0.0   a2 = 0.38689047   ags = 9.179216520e-02 lags = -1.755984120e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.165082675e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.911380500e-10   nfactor = {-7.902623607e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.566332557e-06 wnfactor = 5.273103582e-05 pnfactor = -2.327020611e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.743400046e-03 leta0 = 1.210662561e-9   etab = 4.292802010e-02 letab = -1.897197761e-08 wetab = 1.072026074e-21 petab = -1.767048428e-28   dsub = 1.505414393e+00 ldsub = -2.230393718e-7   voffl = 0.0   minv = 0.0   pclm = 3.786937880e-01 lpclm = 2.637302356e-9   pdiblc1 = 0.39   pdiblc2 = 6.041633520e-03 lpdiblc2 = 1.697666308e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.199682388e-03 lalpha0 = 5.822171861e-10 walpha0 = -5.293955920e-23 palpha0 = -2.524354897e-29   alpha1 = 0.0   beta0 = 1.892222896e+01 lbeta0 = 2.214261161e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.807874800e-01 lkt1 = 6.719886924e-9   kt2 = -4.091695680e-02 lkt2 = 2.864900536e-9   at = 5.149467640e+04 lat = -5.426561953e-4   ute = -1.201588432e+00 lute = 6.927899504e-8   ua1 = 2.302934480e-09 lua1 = 4.477673398e-17   ub1 = -2.697115880e-18 lub1 = 6.311290784e-26   uc1 = -4.599405120e-11 luc1 = 8.798661995e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.22 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.880660082e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.055156887e-07 wvth0 = -6.536389483e-06 pvth0 = 7.928640443e-13   k1 = 4.238027571e-01 lk1 = 3.394183156e-8   k2 = -1.679745637e-01 lk2 = 1.116275303e-08 wk2 = 5.200819131e-07 pk2 = -6.308593606e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.310682975e+05 lvsat = -3.429870278e-02 wvsat = -1.479806403e+00 pvsat = 1.795005167e-7   ua = 6.361200350e-09 lua = -1.060408403e-15 wua = -3.474936317e-14 pua = 4.215097752e-21   ub = -6.228816941e-18 lub = 1.091173308e-24 wub = 4.422776589e-23 pub = -5.364828002e-30   uc = 1.076059409e-10 luc = -8.718430325e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 8.714996960e-02 lu0 = -8.966795562e-09 wu0 = -1.983661761e-07 pu0 = 2.406181716e-14   a0 = 3.952531286e+00 la0 = -4.794420450e-7   keta = 4.955901492e-02 lketa = -1.624955456e-08 pketa = -8.077935669e-28   a1 = 0.0   a2 = 0.38689047   ags = -2.065392429e+00 lags = 3.951095716e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.491611927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.137642643e-9   nfactor = {3.837710627e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.286979768e-06 wnfactor = -1.883251279e-04 pnfactor = 2.284383802e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 6.585351491e-06 lcit = -3.032777402e-13   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.478367509e-01 leta0 = 2.896702053e-08 weta0 = -2.541098842e-21 peta0 = -9.087677628e-28   etab = -1.242688315e-01 letab = 1.301278009e-8   dsub = 3.767858452e-01 ldsub = -7.132730541e-9   voffl = 0.0   minv = 0.0   pclm = 8.348091143e-01 lpclm = -8.461755956e-8   pdiblc1 = -6.670403272e-01 lpdiblc1 = 2.022118146e-7   pdiblc2 = 2.319732429e-02 lpdiblc2 = -1.584217336e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.482554188e-03 lalpha0 = -1.221946710e-10   alpha1 = 0.0   beta0 = 3.068284114e+01 lbeta0 = -3.554394966e-8   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.359701429e-01 lkt1 = -2.098366967e-8   kt2 = -1.682617143e-02 lkt2 = -1.743666706e-9   at = -1.091936143e+04 lat = 1.139714924e-2   ute = 4.592671143e-01 lute = -2.484426710e-7   ua1 = 6.433987771e-09 lua1 = -7.454937607e-16   ub1 = -6.175396171e-18 lub1 = 7.285079276e-25   uc1 = 0.0   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.23 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 5.05e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.907922572e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 8.214148000e-08 wvth0 = 3.672695526e-06 pvth0 = -4.454979673e-13   k1 = 7.630867333e-01 lk1 = -7.213314753e-9   k2 = -2.491551147e-01 lk2 = 2.100995387e-08 wk2 = 3.490450752e-07 pk2 = -4.233916762e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.469883012e+05 lvsat = -1.196979924e-02 wvsat = -2.610115828e-01 pvsat = 3.166070499e-8   ua = 1.481151604e-08 lua = -2.085431696e-15 wua = -8.545367864e-14 pua = 1.036553122e-20   ub = -2.257507078e-17 lub = 3.073973898e-24 wub = 1.257797828e-22 pub = -1.525708766e-29   uc = 8.166707333e-11 luc = -5.572045695e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.179858860e-01 lu0 = -1.270719222e-08 wu0 = -5.268109520e-07 pu0 = 6.390216848e-14   a0 = 0.0   keta = -3.366495898e-02 lketa = -6.154486530e-9   a1 = 0.0   a2 = 0.38689047   ags = 1.009604333e+00 lags = 2.211246437e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.660481612e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.728445837e-9   nfactor = {-2.540630122e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.449947560e-06 wnfactor = 1.417802562e-04 pnfactor = -1.719794508e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.300846521e-06 lcit = 3.377327126e-13   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.811952722e-01 leta0 = -1.094456387e-8   etab = -3.265943586e-02 letab = 1.900560406e-9   dsub = 4.944464162e-01 ldsub = -2.140495780e-8   voffl = 0.0   minv = 0.0   pclm = -2.621870667e-01 lpclm = 4.844807719e-8   pdiblc1 = 1.342867534e+00 lpdiblc1 = -4.159000896e-8   pdiblc2 = 3.207030333e-02 lpdiblc2 = -2.660509694e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.996857262e-03 lalpha0 = -3.058796339e-10   alpha1 = 0.0   beta0 = 3.410467301e+01 lbeta0 = -4.506121549e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.083248333e-01 lkt1 = 1.205295428e-8   kt2 = -8.980038333e-02 lkt2 = 7.108105198e-9   at = 1.090960200e+05 lat = -3.160716526e-3   ute = -2.090441333e+00 lute = 6.083696373e-8   ua1 = -4.245373667e-10 lua1 = 8.644533858e-17   ub1 = 7.279798667e-19 lub1 = -1.088715858e-25   uc1 = 7.856669333e-11 luc1 = -9.530139901e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.24 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.162761188e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.515566545e-8   k1 = 2.427225447e-01 wk1 = 7.898834815e-7   k2 = 5.059433417e-02 wk2 = -3.037806152e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.540631286e+05 wvsat = -5.569378904e-1   ua = -1.514449219e-09 wua = 1.251753307e-15   ub = 2.927791507e-18 wub = -1.341111921e-24   uc = 7.261392233e-11 wuc = -1.089144724e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.116348499e-02 wu0 = 3.790314046e-9   a0 = 2.281552706e+00 wa0 = -1.802539835e-6   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 6.145727805e-01 wags = -2.749062479e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.251289954e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 3.120481283e-8   nfactor = {5.650065209e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.040468635e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.759384422e-05 wcit = -3.806300508e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.313541165e-01 wpclm = 1.001468114e-6   pdiblc1 = 0.39   pdiblc2 = 6.397913279e-03 wpdiblc2 = 9.477688265e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.614451880e-05 walpha0 = 3.832156708e-11   alpha1 = 0.0   beta0 = 1.715499032e+01 wbeta0 = 1.936600023e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.513417791e-01 wkt1 = -1.347430380e-8   kt2 = -3.455331080e-02 wkt2 = -6.851340915e-10   at = -3.121819371e+05 wat = 1.906081105e+0   ute = -1.099546917e+00 wute = -4.879677251e-7   ua1 = 4.201673337e-09 wua1 = -6.397629894e-15   ub1 = -5.071929819e-18 wub1 = 9.016364644e-24   uc1 = 3.160448945e-12 wuc1 = -1.510644546e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.25 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.162761188e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.515566545e-8   k1 = 2.427225447e-01 wk1 = 7.898834815e-7   k2 = 5.059433417e-02 wk2 = -3.037806152e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.540631286e+05 wvsat = -5.569378904e-1   ua = -1.514449219e-09 wua = 1.251753307e-15   ub = 2.927791507e-18 wub = -1.341111921e-24   uc = 7.261392233e-11 wuc = -1.089144724e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.116348499e-02 wu0 = 3.790314046e-9   a0 = 2.281552706e+00 wa0 = -1.802539835e-6   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 6.145727805e-01 wags = -2.749062479e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.251289954e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 3.120481283e-8   nfactor = {5.650065209e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.040468635e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.759384422e-05 wcit = -3.806300508e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = -1.313541165e-01 wpclm = 1.001468114e-6   pdiblc1 = 0.39   pdiblc2 = 6.397913279e-03 wpdiblc2 = 9.477688265e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.614451880e-05 walpha0 = 3.832156708e-11   alpha1 = 0.0   beta0 = 1.715499032e+01 wbeta0 = 1.936600023e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.513417791e-01 wkt1 = -1.347430380e-8   kt2 = -3.455331080e-02 wkt2 = -6.851340915e-10   at = -3.121819371e+05 wat = 1.906081105e+0   ute = -1.099546917e+00 wute = -4.879677251e-7   ua1 = 4.201673337e-09 wua1 = -6.397629894e-15   ub1 = -5.071929819e-18 wub1 = 9.016364644e-24   uc1 = 3.160448945e-12 wuc1 = -1.510644546e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.26 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.156394467e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.509316099e-09 wvth0 = 3.502732852e-08 pvth0 = 3.991881435e-14   k1 = -8.028418694e-02 lk1 = 1.273066432e-06 wk1 = 1.946806013e-06 pk1 = -4.559778772e-12   k2 = 1.695112125e-01 lk2 = -4.686870924e-07 wk2 = -7.420164709e-07 pk2 = 1.727218978e-12   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.350619352e+05 lvsat = -1.107500596e+00 wvsat = -1.019921189e+00 pvsat = 1.824756074e-6   ua = -1.747066623e-09 lua = 9.168149766e-16 wua = 2.349875105e-15 pua = -4.328027441e-21   ub = 3.060098871e-18 lub = -5.214630113e-25 wub = -2.102122661e-24 pub = 2.999371627e-30   uc = 3.868671549e-11 luc = 1.337173003e-16 wuc = 3.326097123e-17 puc = -1.740179269e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.891256240e-02 lu0 = 8.871561231e-09 wu0 = 1.264755097e-08 pu0 = -3.490902790e-14   a0 = 2.520441035e+00 la0 = -9.415305700e-07 wa0 = -3.021968843e-06 pa0 = 4.806135549e-12   keta = 1.568695494e-01 lketa = -6.182699552e-07 wketa = 2.646062198e-07 pketa = -1.042892494e-12   a1 = 0.0   a2 = 0.38689047   ags = 3.854502911e-01 lags = 9.030404675e-07 wags = -3.308186878e-06 pags = 1.195506895e-11   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.481622661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.078102982e-08 wvoff = 1.099094612e-07 pvoff = -3.101986308e-13   nfactor = {-4.030135264e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.815257413e-06 wnfactor = 4.823713752e-06 pnfactor = -1.096960398e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 2.981805911e-05 lcit = -4.817929816e-11 wcit = -7.500886096e-11 pcit = 1.456147018e-16   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374486321e-01 letab = 2.658352936e-07 wetab = -5.785721031e-11 petab = 2.280326230e-16   dsub = 5.808742267e-01 ldsub = -8.227158985e-08 wdsub = 5.699045314e-07 pdsub = -2.246164730e-12   voffl = 0.0   minv = 0.0   pclm = -1.085007159e-01 lpclm = -9.007210793e-08 wpclm = 9.800395177e-07 ppclm = 8.445652704e-14   pdiblc1 = 0.39   pdiblc2 = 2.902643952e-03 lpdiblc2 = 1.377590500e-08 wpdiblc2 = 7.781274331e-09 ppdiblc2 = -2.693289524e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.475066708e-05 lalpha0 = 3.188321961e-10 walpha0 = -1.990092691e-11 palpha0 = 2.294723156e-16   alpha1 = 0.0   beta0 = 1.333870485e+01 lbeta0 = 1.504112590e-05 wbeta0 = 2.693783172e-06 pbeta0 = -2.984285944e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.220501773e-01 lkt1 = -1.154469904e-07 wkt1 = -1.088685037e-07 pkt1 = 3.759771600e-13   kt2 = -6.811115124e-02 lkt2 = 1.322615165e-07 wkt2 = 1.050391271e-07 pkt2 = -4.166910306e-13   at = -6.945766975e+05 lat = 1.507132469e+00 wat = 3.870773051e+00 pat = -7.743440366e-6   ute = -9.355685643e-01 lute = -6.462878816e-07 wute = -1.132303452e-06 pute = 2.539520399e-12   ua1 = 5.136454936e-09 lua1 = -3.684254719e-15 wua1 = -9.644431709e-15 pua1 = 1.279661999e-20   ub1 = -6.649892702e-18 lub1 = 6.219225109e-24 wub1 = 1.499124846e-23 pub1 = -2.354880957e-29   uc1 = 2.394830587e-11 luc1 = -8.193118050e-17 wuc1 = -1.943428301e-16 puc1 = 1.705730617e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.27 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.100884862e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.328539564e-08 wvth0 = 7.331070604e-08 pvth0 = -3.440070644e-14   k1 = 7.102349569e-01 lk1 = -2.615683823e-07 wk1 = -7.957072887e-07 pk1 = 7.642622999e-13   k2 = -1.175636857e-01 lk2 = 8.861140740e-08 wk2 = 2.947329214e-07 pk2 = -2.854226171e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.163652801e+04 lvsat = 5.690146675e-03 wvsat = -1.849905850e-01 pvsat = 2.039052929e-7   ua = -9.730026545e-10 lua = -5.858754064e-16 wua = -7.321245649e-17 pua = 3.759124419e-22   ub = 2.766016797e-18 lub = 4.943851763e-26 wub = -7.900483932e-25 pub = 4.522418524e-31   uc = 1.333320618e-10 luc = -5.001771041e-17 wuc = -9.046635467e-17 puc = 6.617393085e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.773892243e-02 lu0 = -8.263051495e-09 wu0 = -8.528571555e-09 pu0 = 6.200178762e-15   a0 = 1.977844788e+00 la0 = 1.118115254e-07 wa0 = 5.007015098e-07 pa0 = -2.032424407e-12   keta = -1.779157995e-01 lketa = 3.164884269e-08 wketa = -4.121242262e-07 pketa = 2.708443207e-13   a1 = 0.0   a2 = 0.38689047   ags = -1.774618494e-01 lags = 1.995821806e-06 wags = 5.179170437e-06 pags = -4.521437809e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.885902271e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.434435652e-08 wvoff = -9.290929682e-08 pvoff = 8.353342423e-14   nfactor = {1.667426061e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.040869584e-07 wnfactor = -2.525568453e-06 pnfactor = 3.297557565e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.161082290e-04 leta0 = -3.127090491e-11 weta0 = 4.858372626e-11 peta0 = -9.431558779e-17   etab = -5.402721130e-04 letab = 5.509439083e-11 wetab = 9.013272405e-11 petab = -5.926023658e-17   dsub = -2.029035086e-01 ldsub = 1.439276128e-06 wdsub = 3.988974535e-07 pdsub = -1.914188689e-12   voffl = 0.0   minv = 0.0   pclm = -8.201668524e-01 lpclm = 1.291485363e-06 wpclm = 3.300845917e-06 ppclm = -4.420924936e-12   pdiblc1 = 0.39   pdiblc2 = 9.806762754e-03 lpdiblc2 = 3.729391665e-10 wpdiblc2 = -2.043316273e-08 ppdiblc2 = 2.783979142e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.383292683e-04 lalpha0 = -5.599388256e-11 walpha0 = 2.806660507e-10 palpha0 = -3.540183580e-16   alpha1 = 0.0   beta0 = 2.034207087e+01 lbeta0 = 1.445491455e-06 wbeta0 = 5.275984448e-06 pbeta0 = -7.997113283e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.987152587e-01 lkt1 = 3.338293223e-08 wkt1 = 1.701483546e-07 pkt1 = -1.656782671e-13   kt2 = 5.456549607e-02 lkt2 = -1.058906589e-07 wkt2 = -3.179859875e-07 pkt2 = 4.045276243e-13   at = 9.415439160e+04 lat = -2.403119392e-02 wat = -2.533145157e-01 pat = 2.626508279e-7   ute = -1.263480958e+00 lute = -9.711552635e-09 wute = -1.351420905e-07 pute = 6.037310487e-13   ua1 = 4.986475602e-09 lua1 = -3.393099838e-15 wua1 = -9.675231151e-15 pua1 = 1.285641095e-20   ub1 = -5.944652660e-18 lub1 = 4.850142615e-24 wub1 = 1.200501798e-23 pub1 = -1.775164035e-29   uc1 = -9.437225678e-11 luc1 = 1.477645278e-16 wuc1 = 2.212620611e-16 puc1 = -6.362407137e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.28 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.259748119e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.668402709e-09 wvth0 = 6.747985084e-08 pvth0 = -2.891212244e-14   k1 = 4.045527039e-01 lk1 = 2.617032237e-08 wk1 = 1.184090302e-07 pk1 = -9.619539105e-14   k2 = -1.289021520e-03 lk2 = -2.083793400e-08 wk2 = -7.625099717e-08 pk2 = 6.378454547e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -5.132826550e+04 lvsat = 1.120239068e-01 wvsat = 1.921834095e-01 pvsat = -1.511285881e-7   ua = -1.092645942e-09 lua = -4.732551794e-16 wua = -1.814574561e-15 pua = 2.015056591e-21   ub = 2.593696377e-18 lub = 2.116437294e-25 wub = 1.646597911e-24 pub = -1.841373314e-30   uc = 9.168043527e-11 luc = -1.081103439e-17 wuc = 1.224750255e-17 puc = -3.051062295e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.556077116e-02 lu0 = -6.212757709e-09 wu0 = -1.857534552e-08 pu0 = 1.565720709e-14   a0 = 2.889210684e+00 la0 = -7.460571934e-07 wa0 = -4.743494296e-06 pa0 = 2.903937105e-12   keta = -2.878701494e-01 lketa = 1.351488722e-07 wketa = -1.528583128e-07 pketa = 2.679731642e-14   a1 = 0.0   a2 = 0.38689047   ags = 4.625262814e+00 lags = -2.524982920e-06 wags = -4.373112187e-06 pags = 4.470125826e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.104352106e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.034690842e-09 wvoff = -3.035755363e-08 pvoff = 2.465346837e-14   nfactor = {6.331202753e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.695050776e-07 wnfactor = 1.539701833e-06 pnfactor = -5.290813547e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 9.224882881e-04 leta0 = -4.137963677e-10 weta0 = -1.643562691e-10 peta0 = 1.061248298e-16   etab = -8.999025590e-04 letab = 3.936145297e-10 wetab = 2.950630436e-10 petab = -2.521611464e-16   dsub = 1.613966110e+00 ldsub = -2.709432444e-07 wdsub = -3.077413033e-06 pdsub = 1.358062371e-12   voffl = 0.0   minv = 0.0   pclm = 5.780759410e-01 lpclm = -2.468057857e-08 wpclm = -2.019484181e-06 ppclm = 5.871017851e-13   pdiblc1 = 0.39   pdiblc2 = 1.185760567e-02 lpdiblc2 = -1.557519268e-09 wpdiblc2 = 1.030913168e-08 ppdiblc2 = -1.097930302e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.943817368e-05 lalpha0 = 4.650530485e-11 walpha0 = -1.124991166e-10 palpha0 = 1.606801390e-17   alpha1 = 0.0   beta0 = 1.979734008e+01 lbeta0 = 1.958246545e-06 wbeta0 = -4.756723766e-06 pbeta0 = 1.446674960e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.515876842e-01 lkt1 = -1.097825368e-08 wkt1 = -5.927681196e-08 pkt1 = 5.027964226e-14   kt2 = -6.593436738e-02 lkt2 = 7.535862564e-09 wkt2 = 1.465652962e-07 pkt2 = -3.275449903e-14   at = 1.137774712e+05 lat = -4.250239872e-02 wat = -9.668921979e-02 pat = 1.152194368e-7   ute = -2.143238017e+00 lute = 8.184037670e-07 wute = 4.297030998e-06 pute = -3.568273480e-12   ua1 = -2.348402038e-09 lua1 = 3.511220485e-15 wua1 = 2.167124227e-14 pua1 = -1.665002448e-20   ub1 = 4.098342711e-18 lub1 = -4.603328927e-24 wub1 = -2.961988330e-23 pub1 = 2.142987923e-29   uc1 = 1.757880365e-10 luc1 = -1.065373563e-16 wuc1 = -1.031000652e-15 puc1 = 5.425141778e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.29 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.937468020e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.157618198e-08 wvth0 = 1.601900722e-09 pvth0 = 1.598169451e-16   k1 = 3.459336161e-01 lk1 = 5.203892582e-08 wk1 = -1.115932767e-07 pk1 = 5.304626971e-15   k2 = -2.391408515e-02 lk2 = -1.085349342e-08 wk2 = 8.604124844e-08 pk2 = -7.835022518e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.501438671e+05 lvsat = -2.101574530e-02 wvsat = -2.785377236e-01 pvsat = 5.660064793e-8   ua = -3.008159957e-09 lua = 3.720611554e-16 wua = 7.371401141e-15 pua = -2.038714487e-21   ub = 3.691302112e-18 lub = -2.727296816e-25 wub = -6.140006870e-24 pub = 1.594855376e-30   uc = 5.424176768e-11 luc = 5.710649622e-18 wuc = -1.580443455e-17 puc = -1.813130311e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.223402730e-02 lu0 = 4.081334356e-09 wu0 = 5.965296638e-08 pu0 = -1.886494695e-14   a0 = 1.065157185e+00 la0 = 5.889761606e-08 wa0 = 2.961539856e-06 pa0 = -4.962944667e-13   keta = 6.202044834e-02 lketa = -1.925784853e-08 wketa = -1.751555097e-07 pketa = 3.663706938e-14   a1 = 0.0   a2 = 0.38689047   ags = -1.935417760e+00 lags = 3.702454175e-07 wags = 1.016108567e-05 pags = -1.943815689e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.241608290e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.022424557e-09 wvoff = 3.835731673e-08 pvoff = -5.670403924e-15   nfactor = {2.689695783e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.380616940e-07 wnfactor = -3.613762749e-07 pnfactor = 3.098644142e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.600656514e-03 leta0 = -1.154371932e-09 weta0 = -2.678628197e-08 peta0 = 1.185438064e-14   etab = 8.676520821e-02 letab = -3.829299885e-08 wetab = -2.197273298e-07 petab = 9.684372082e-14   dsub = 1.417871537e+00 ldsub = -1.844067092e-07 wdsub = 4.387954372e-07 pdsub = -1.936404265e-13   voffl = 0.0   minv = 0.0   pclm = 5.863177459e-01 lpclm = -2.831768708e-08 wpclm = -1.040683945e-06 ppclm = 1.551572413e-13   pdiblc1 = 0.39   pdiblc2 = 5.821920400e-03 lpdiblc2 = 1.106028641e-09 wpdiblc2 = 1.101279058e-09 ppdiblc2 = 2.965495059e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -9.800230863e-04 lalpha0 = 4.919805589e-10 walpha0 = -1.101009301e-09 palpha0 = 4.522975583e-16   alpha1 = 0.0   beta0 = 1.941145577e+01 lbeta0 = 2.128537294e-06 wbeta0 = -2.452175985e-06 pbeta0 = 4.296780237e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.294973675e-01 lkt1 = 2.340328958e-08 wkt1 = 2.441510048e-07 pkt1 = -8.362305329e-14   kt2 = -5.783219499e-02 lkt2 = 3.960373886e-09 wkt2 = 8.478509413e-08 pkt2 = -5.490895845e-15   at = 2.583131587e+03 lat = 6.567663337e-03 wat = 2.451617816e-01 pat = -3.563941011e-8   ute = -8.577533084e-01 lute = 2.511193653e-07 wute = -1.723421982e-06 pute = -9.114475799e-13   ua1 = 5.024960738e-09 lua1 = 2.573554915e-16 wua1 = -1.364374832e-14 pua1 = -1.065519135e-21   ub1 = -6.543737276e-18 lub1 = 9.302097145e-26 wub1 = 1.928061275e-23 pub1 = -1.499096826e-31   uc1 = -1.508887272e-10 luc1 = 3.762509953e-17 wuc1 = 5.257688293e-16 puc1 = -1.444881942e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.30 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.161226294e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.498667775e-08 wvth0 = -1.980851832e-07 pvth0 = 3.835995611e-14   k1 = 4.399985349e-01 lk1 = 3.404430685e-08 wk1 = -8.117890650e-08 pk1 = -5.136420489e-16   k2 = -7.646866175e-02 lk2 = -7.998029160e-10 wk2 = 6.142230558e-08 pk2 = -3.125418749e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.079825995e+05 lvsat = 6.179705195e-03 wvsat = 1.396121951e-01 pvsat = -2.339143152e-8   ua = 1.678023323e-09 lua = -5.244057062e-16 wua = -1.127564080e-14 pua = 1.528464636e-21   ub = 1.133386590e-18 lub = 2.165995579e-25 wub = 7.325825020e-24 pub = -9.811582645e-31   uc = 1.764838944e-10 luc = -1.767426922e-17 wuc = -3.452404105e-16 puc = 4.488979910e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.225729567e-02 lu0 = -7.401116883e-09 wu0 = -1.237188819e-07 pu0 = 1.621408763e-14   a0 = 3.752316936e+00 la0 = -4.551560443e-07 wa0 = 1.003544398e-06 pa0 = -1.217299354e-13   keta = -2.930997983e-02 lketa = -1.786337623e-09 wketa = 3.953190058e-07 pketa = -7.249470544e-14   a1 = 0.0   a2 = 0.38689047   ags = -2.198035624e+00 lags = 4.204842149e-07 wags = 6.648541224e-07 pags = -1.271865936e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.594343399e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.770247196e-09 wvoff = 5.149260951e-08 pvoff = -8.183185433e-15   nfactor = {-5.153086073e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.750556459e-07 wnfactor = 6.617267758e-06 pnfactor = -1.025150189e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 8.993133942e-06 lcit = -7.638865232e-13 wcit = -1.206864837e-11 pcit = 2.308732433e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.954175230e-01 leta0 = 3.672650577e-08 weta0 = 2.384914830e-07 peta0 = -3.889325580e-14   etab = -2.747495643e-01 letab = 3.086477713e-08 wetab = 7.542621013e-07 petab = -8.948045735e-14   dsub = 7.353697166e-01 ldsub = -5.384411098e-08 wdsub = -1.797347867e-06 pdsub = 2.341337877e-13   voffl = 0.0   minv = 0.0   pclm = 1.154913403e+00 lpclm = -1.370900363e-07 wpclm = -1.604474732e-06 ppclm = 2.630104187e-13   pdiblc1 = -6.748561169e-01 lpdiblc1 = 2.037069752e-07 wpdiblc1 = 3.917547384e-08 ppdiblc1 = -7.494268145e-15   pdiblc2 = 1.987436220e-02 lpdiblc2 = -1.582203475e-09 wpdiblc2 = 1.665584902e-08 ppdiblc2 = -1.009417410e-17   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.549111578e-04 lalpha0 = 4.297866470e-10 walpha0 = 1.572607443e-08 palpha0 = -2.766723559e-15   alpha1 = 0.0   beta0 = 2.621406602e+01 lbeta0 = 8.271979521e-07 wbeta0 = 2.239906497e-05 pbeta0 = -4.324364371e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.367254008e-02 lkt1 = -3.701399992e-08 wkt1 = -6.129983893e-07 pkt1 = 8.034962580e-14   kt2 = -2.275921805e-02 lkt2 = -2.749086602e-09 wkt2 = 2.973850624e-08 pkt2 = 5.039516417e-15   at = -7.615927262e+04 lat = 2.163108526e-02 wat = 3.270052689e-01 pat = -5.129606921e-8   ute = 3.641871050e+00 lute = -6.096587745e-07 wute = -1.595232484e-05 pute = 1.810541537e-12   ua1 = 1.608591655e-08 lua1 = -1.858605355e-15 wua1 = -4.837884521e-14 pua1 = 5.579304901e-21   ub1 = -1.520665470e-17 lub1 = 1.750237074e-24 wub1 = 4.526782866e-23 pub1 = -5.121264086e-30   uc1 = 1.094121817e-10 luc1 = -1.217046436e-17 wuc1 = -5.484121491e-16 puc1 = 6.100262702e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.31 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.01e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {1.578560245e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.010614271e-10 wvth0 = 4.214433110e-07 pvth0 = -3.678885025e-14   k1 = 6.662845079e-01 lk1 = 6.595818329e-09 wk1 = 4.852066348e-07 pk1 = -6.921620820e-14   k2 = -1.744377166e-01 lk2 = 1.108384344e-08 wk2 = -2.546467534e-08 pk2 = 7.413972037e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.366499493e+05 lvsat = -9.427644332e-03 wvsat = -2.091921444e-01 pvsat = 1.891853486e-8   ua = -3.087045757e-09 lua = 5.359717327e-17 wua = 4.260177582e-15 pua = -3.560301333e-22   ub = 1.900468845e-18 lub = 1.235524803e-25 wub = 3.099811827e-24 pub = -4.685428642e-31   uc = 9.475204280e-11 luc = -7.760195622e-18 wuc = -6.558644670e-17 puc = 1.096777328e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -4.359501379e-03 lu0 = 1.892500599e-09 wu0 = 8.642695048e-08 pu0 = -9.276601838e-15   a0 = 0.0   keta = -2.163792710e-01 lketa = 2.090516740e-08 wketa = 9.158280821e-07 pketa = -1.356324564e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.298767796e+00 lags = -3.678039968e-09 wags = -1.449388483e-06 pags = 1.292710344e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {1.198147239e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.510266425e-08 wvoff = -7.339059815e-07 pvoff = 8.708566366e-14   nfactor = {5.740314171e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.837513971e-07 wnfactor = -1.433748145e-05 pnfactor = 1.516660889e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.879328671e-05 lcit = -1.952645054e-12 wcit = -8.767823260e-11 pcit = 1.148017500e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.298200805e-01 leta0 = -2.698481554e-08 weta0 = -7.449595579e-07 peta0 = 8.039935546e-14   etab = 8.702131265e-03 letab = -3.517913544e-09 wetab = -2.073186510e-07 petab = 2.715928790e-14   dsub = 3.872745213e-01 ldsub = -1.162016380e-08 wdsub = 5.371830471e-07 pdsub = -4.904481220e-14   voffl = 0.0   minv = 0.0   pclm = -1.181273222e+00 lpclm = 1.462894013e-07 wpclm = 4.606781491e-06 ppclm = -4.904149612e-13   pdiblc1 = 1.881849870e+00 lpdiblc1 = -1.064214611e-07 wpdiblc1 = -2.701568115e-06 ppdiblc1 = 3.249579292e-13   pdiblc2 = 3.212283805e-02 lpdiblc2 = -3.067943597e-09 wpdiblc2 = -2.633224067e-10 ppdiblc2 = 2.042201320e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 8.267147417e-03 lalpha0 = -6.524590581e-10 walpha0 = -2.140418886e-08 palpha0 = 1.737177377e-15   alpha1 = 0.0   beta0 = 3.922057217e+01 lbeta0 = -7.504912441e-07 wbeta0 = -2.564267719e-05 pbeta0 = 1.503098953e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -8.154066230e-01 lkt1 = 6.023634434e-08 wkt1 = 2.040436408e-06 pkt1 = -2.415120151e-13   kt2 = -1.459355176e-01 lkt2 = 1.219219853e-08 wkt2 = 2.813689402e-07 pkt2 = -2.548325522e-14   at = 2.447254444e+05 lat = -1.729223091e-02 wat = -6.798221454e-01 pat = 7.083209613e-8   ute = -2.368722817e+00 lute = 1.194262616e-07 wute = 1.394844197e-06 pute = -2.936700673e-13   ua1 = -2.092406846e-10 lua1 = 1.179972173e-16 wua1 = -1.079142324e-15 pua1 = -1.581490594e-22   ub1 = 4.872247405e-20 lub1 = -1.002401768e-25 wub1 = 3.404675792e-24 pub1 = -4.326364293e-32   uc1 = 5.337504057e-11 luc1 = -5.373159133e-18 wuc1 = 1.262693807e-16 puc1 = -2.083624255e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.32 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4312167+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.50407   k2 = -0.049917061   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169790.0   ua = -1.10028365e-9   ub = 2.48406e-18   uc = 6.9010287e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03241758   a0 = 1.6851493   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.523615   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.24013304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0067115   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.8823913e-5   alpha1 = 0.0   beta0 = 17.79575   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.2558   kt2 = -0.03478   at = 318480.0   ute = -1.261   ua1 = 2.0849e-9   ub1 = -2.0887e-18   uc1 = -4.6822e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.33 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4312167+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.50407   k2 = -0.049917061   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169790.0   ua = -1.10028365e-9   ub = 2.48406e-18   uc = 6.9010287e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03241758   a0 = 1.6851493   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.523615   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.24013304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0067115   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.8823913e-5   alpha1 = 0.0   beta0 = 17.79575   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.2558   kt2 = -0.03478   at = 318480.0   ute = -1.261   ua1 = 2.0849e-9   ub1 = -2.0887e-18   uc1 = -4.6822e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.34 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.272288815e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.571718890e-8   k1 = 5.638523335e-01 lk1 = -2.356201110e-7   k2 = -7.599856336e-02 lk2 = 1.027950253e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.976022800e+05 lvsat = -5.037465394e-1   ua = -9.695672919e-10 lua = -5.151923821e-16   ub = 2.364572985e-18 lub = 4.709341722e-25   uc = 4.969171863e-11 luc = 7.614027353e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.309723690e-02 lu0 = -2.678731721e-9   a0 = 1.520567148e+00 la0 = 6.486676363e-7   keta = 2.444193765e-01 lketa = -9.633300886e-7   a1 = 0.0   a2 = 0.38689047   ags = -7.091240891e-01 lags = 4.858594572e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.117967024e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.185388367e-8   nfactor = {1.193000751e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.857624900e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374677752e-01 letab = 2.659107424e-7   dsub = 7.694376067e-01 ldsub = -8.254564393e-7   voffl = 0.0   minv = 0.0   pclm = 2.157633560e-01 lpclm = -6.212811500e-8   pdiblc1 = 0.39   pdiblc2 = 5.477221460e-03 lpdiblc2 = 4.864662010e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -6.133525421e-05 lalpha0 = 3.947573257e-10 palpha0 = 2.524354897e-29   alpha1 = 0.0   beta0 = 1.422999248e+01 lbeta0 = 1.405372009e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.580713210e-01 lkt1 = 8.951957457e-9   kt2 = -3.335702710e-02 lkt2 = -5.608363091e-9   at = 5.861396494e+05 lat = -1.054926976e+0   ute = -1.310211955e+00 lute = 1.939590782e-7   ua1 = 1.945417595e-09 lua1 = 5.497420028e-16   ub1 = -1.689762850e-18 lub1 = -1.572330989e-24   uc1 = -4.035358840e-11 luc1 = -2.549395064e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.35 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.343446796e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.903290177e-9   k1 = 4.469605880e-01 lk1 = -8.698165484e-9   k2 = -2.004588617e-02 lk2 = -5.825906982e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.289958000e+02 lvsat = 7.315595735e-2   ua = -9.972263402e-10 lua = -4.614978717e-16   ub = 2.504614778e-18 lub = 1.990710395e-25   uc = 1.033996070e-10 luc = -2.812285017e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.491708791e-02 lu0 = -6.211608491e-9   a0 = 2.143511077e+00 la0 = -5.606534132e-7   keta = -3.142746680e-01 lketa = 1.212626600e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.536161800e+00 lags = 4.998210752e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.195997697e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.294210896e-9   nfactor = {8.317953586e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.869705185e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.321830470e-04 leta0 = -6.247694914e-11 weta0 = -1.058791184e-22   etab = -5.104500460e-04 letab = 3.548705330e-11   dsub = -7.092096076e-02 ldsub = 8.059316477e-7   voffl = 0.0   minv = 0.0   pclm = 2.719786360e-01 lpclm = -1.712588381e-7   pdiblc1 = 0.39   pdiblc2 = 3.046075630e-03 lpdiblc2 = 9.584245409e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.311927854e-04 lalpha0 = -1.731273575e-10   alpha1 = 0.0   beta0 = 2.208772721e+01 lbeta0 = -1.200500334e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.424185510e-01 lkt1 = -2.143476494e-8   kt2 = -5.064600740e-02 lkt2 = 2.795473437e-8   at = 1.034063220e+04 lat = 6.287165581e-2   ute = -1.308195200e+00 lute = 1.900439518e-7   ua1 = 1.785247700e-09 lua1 = 8.606798200e-16   ub1 = -1.972572000e-18 lub1 = -1.023313586e-24   uc1 = -2.116364060e-11 luc1 = -6.274739630e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.36 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.483017597e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.123450936e-8   k1 = 4.437305060e-01 lk1 = -5.657689298e-9   k2 = -2.651806421e-02 lk2 = 2.663542088e-10   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.225914480e+04 lvsat = 6.202023810e-2   ua = -1.693031259e-09 lua = 1.934632981e-16   ub = 3.138503534e-18 lub = -3.976084466e-25   uc = 9.573274640e-11 luc = -2.090603429e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.941477698e-02 lu0 = -1.032283213e-9   a0 = 1.319738487e+00 la0 = 2.147637257e-7   keta = -3.384461293e-01 lketa = 1.440152565e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.178338339e+00 lags = -1.045959701e-06 wags = 4.336808690e-19   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.204795647e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.122361904e-9   nfactor = {1.142558902e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.944487953e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.681079060e-04 leta0 = -3.786830189e-10   etab = -8.022755325e-04 letab = 3.101823837e-10   dsub = 5.957474947e-01 ldsub = 1.783966306e-7   voffl = 0.0   minv = 0.0   pclm = -9.010748600e-02 lpclm = 1.695728286e-07 ppclm = 1.292469707e-26   pdiblc1 = 0.39   pdiblc2 = 1.526857120e-02 lpdiblc2 = -1.920789671e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -7.784224971e-06 lalpha0 = 5.182170233e-11   alpha1 = 0.0   beta0 = 1.822349067e+01 lbeta0 = 2.436905523e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.712005060e-01 lkt1 = 5.657689298e-9   kt2 = -1.744054760e-02 lkt2 = -3.301564944e-9   at = 8.178606720e+04 lat = -4.379932155e-3   ute = -7.214864000e-01 lute = -3.622250417e-7   ua1 = 4.821926438e-09 lua1 = -1.997745876e-15 pua1 = -3.851859889e-34   ub1 = -5.701939620e-18 lub1 = 2.487140154e-24   uc1 = -1.653374624e-10 luc1 = 7.296342216e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.37 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.942768203e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.152330361e-8   k1 = 3.090109312e-01 lk1 = 5.379405906e-8   k2 = 4.554241956e-03 lk2 = -1.344585450e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.579845461e+05 lvsat = -2.288381513e-3   ua = -5.691965212e-10 lua = -3.024849716e-16   ub = 1.659768084e-18 lub = 2.549575076e-25   uc = 4.901258028e-11 luc = -2.884249758e-19   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.197130670e-02 lu0 = -2.160479778e-9   a0 = 2.045037032e+00 la0 = -1.053105222e-7   keta = 4.067031414e-03 lketa = -7.135801324e-9   a1 = 0.0   a2 = 0.38689047   ags = 1.426564032e+00 lags = -2.729016993e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.114696064e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.462672875e-10   nfactor = {2.570127806e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.553736221e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -6.262077039e-03 leta0 = 2.767867597e-09 weta0 = -5.293955920e-23 peta0 = -7.967495143e-29   etab = 1.406438606e-02 letab = -6.250475379e-09 wetab = 2.646977960e-22 petab = -4.038967835e-28   dsub = 1.563055065e+00 ldsub = -2.484762003e-7   voffl = 0.0   minv = 0.0   pclm = 2.419883514e-01 lpclm = 2.301893551e-8   pdiblc1 = 0.39   pdiblc2 = 6.186298800e-03 lpdiblc2 = 2.087217140e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.344312232e-03 lalpha0 = 6.416315120e-10 palpha0 = 4.417621069e-29   alpha1 = 0.0   beta0 = 1.860010831e+01 lbeta0 = 2.270704159e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.487155240e-01 lkt1 = -4.264933259e-9   kt2 = -2.977948960e-02 lkt2 = 2.143610160e-9   at = 8.369940920e+04 lat = -5.224289980e-3   ute = -1.427979120e+00 lute = -5.044980434e-8   ua1 = 5.106760540e-10 lua1 = -9.519108163e-17   ub1 = -1.643924768e-19 lub1 = 4.342060001e-26   uc1 = 2.307154520e-11 luc1 = -1.018147290e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.38 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.505825089e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.229458183e-8   k1 = 4.131390029e-01 lk1 = 3.387435895e-8   k2 = -5.614596399e-02 lk2 = -1.833905104e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.541758581e+05 lvsat = -1.559779482e-3   ua = -2.052729501e-09 lua = -1.868511253e-17   ub = 3.557270329e-18 lub = -1.080346719e-25   uc = 6.225476458e-11 luc = -2.821654834e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.132263161e-02 lu0 = -2.036388235e-9   a0 = 4.084358029e+00 la0 = -4.954326289e-7   keta = 1.014885729e-01 lketa = -2.577254221e-8   a1 = 0.0   a2 = 0.38689047   ags = -1.978056429e+00 lags = 3.784021948e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.423970645e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.062690019e-9   nfactor = {1.674135950e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.358658799e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.165082362e-01 leta0 = 2.385795785e-08 weta0 = 3.388131789e-21 peta0 = -8.077935669e-28   etab = -2.518809681e-02 letab = 1.258524594e-9   dsub = 1.406841681e-01 ldsub = 2.362335233e-8   voffl = 0.0   minv = 0.0   pclm = 6.240434735e-01 lpclm = -5.006820933e-8   pdiblc1 = -6.618941920e-01 lpdiblc1 = 2.012273589e-7   pdiblc2 = 2.538525571e-02 lpdiblc2 = -1.585543318e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.548349361e-03 lalpha0 = -4.856346507e-10   alpha1 = 0.0   beta0 = 3.362520800e+01 lbeta0 = -6.035974128e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.164943143e-01 lkt1 = -1.042885068e-8   kt2 = -1.291968714e-02 lkt2 = -1.081670050e-9   at = 3.203642571e+04 lat = 4.658838761e-3   ute = -1.636248571e+00 lute = -1.060785829e-8   ua1 = 7.888718143e-11 lua1 = -1.258987031e-17 pua1 = 7.523163845e-37   ub1 = -2.289622829e-19 lub1 = 5.577280391e-26 pub1 = 2.802596929e-45   uc1 = -7.204004886e-11 luc1 = 8.013375046e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.39 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 3.01e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-5.322431424e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.701020082e-07 wvth0 = 1.698479008e-05 pvth0 = -2.060255037e-12   k1 = 8.268240333e-01 lk1 = -1.630563524e-8   k2 = 1.561728285e+00 lk2 = -1.980820515e-07 wk2 = -5.272765991e-06 pk2 = 6.395865147e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.618663619e+06 lvsat = -1.792021448e-01 wvsat = -4.386121158e+00 pvsat = 5.320364964e-7   ua = 8.172397655e-08 lua = -1.018079956e-14 wua = -2.520684157e-13 pua = 3.057589882e-20   ub = -9.516889629e-17 lub = 1.186744934e-23 wub = 2.964774075e-22 pub = -3.596270953e-29   uc = 7.305156248e-11 luc = -4.131306418e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.834040750e-01 lu0 = -3.261386732e-08 wu0 = -7.832952946e-07 pu0 = 9.501371923e-14   a0 = 0.0   keta = 8.663926820e-02 lketa = -2.397132155e-8   a1 = 0.0   a2 = 0.38689047   ags = 8.192110000e-01 lags = 3.909365570e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.230115475e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.711226815e-9   nfactor = {1.719719585e+02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.052126000e-05 wnfactor = -5.167476917e-04 pnfactor = 6.268149500e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.021666667e-05 lcit = 1.845781667e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 8.333653029e-02 leta0 = -3.832123299e-10   etab = -5.989305161e-02 letab = 5.468235612e-9   dsub = 5.650113973e-01 ldsub = -2.784754057e-8   voffl = 0.0   minv = 0.0   pclm = 3.429650333e-01 lpclm = -1.597339454e-8   pdiblc1 = 9.879864480e-01 lpdiblc1 = 1.096837298e-9   pdiblc2 = 3.203571300e-02 lpdiblc2 = -2.392243787e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.185178467e-03 lalpha0 = -7.768202129e-11   alpha1 = 0.0   beta0 = 3.073622152e+01 lbeta0 = -2.531633527e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.402907667e-01 lkt1 = -1.967234100e-8   kt2 = -5.283943667e-02 lkt2 = 3.760595568e-9   at = 1.979380333e+04 lat = 6.143868856e-3   ute = -1.907213000e+00 lute = 2.226012690e-8   ua1 = -5.662947400e-10 lua1 = 6.567069676e-17 wua1 = -2.524354897e-29 pua1 = -3.009265538e-36   ub1 = 1.175221983e-18 lub1 = -1.145547476e-25   uc1 = 9.515358400e-11 luc1 = -1.226721262e-17 wuc1 = -3.155443621e-30 puc1 = -3.761581923e-37   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.40 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.412257709e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -3.015082478e-8   k1 = 4.681262989e-01 wk1 = 1.082750080e-7   k2 = -4.122919261e-02 wk2 = -2.617090033e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.319130474e+05 wvsat = 1.140986381e-1   ua = -1.249558358e-09 wua = 4.496676663e-16   ub = 2.609314994e-18 wub = -3.773118814e-25   uc = 1.264656591e-10 wuc = -1.730756901e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.260217473e-02 wu0 = -5.560639416e-10   a0 = 1.387952274e+00 wa0 = 8.952614623e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.672929384e-01 wags = -1.315732378e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.204319435e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.695240176e-8   nfactor = {8.491646233e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.177733710e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.156851852e-06 wcit = 1.854659268e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 5.655476770e-03 wpdiblc2 = 3.181111576e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.523936430e-05 walpha0 = 1.079791528e-11   alpha1 = 0.0   beta0 = 1.779868928e+01 wbeta0 = -8.854143344e-9   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.535465922e-01 wkt1 = -6.788052919e-9   kt2 = -3.282950933e-02 wkt2 = -5.875560560e-9   at = 6.389441389e+05 wat = -9.653501488e-1   ute = -1.359755904e+00 wute = 2.974873465e-7   ua1 = 2.234265226e-09 wua1 = -4.499403383e-16   ub1 = -2.855474330e-18 wub1 = 2.309792652e-24   uc1 = -1.825682696e-10 wuc1 = 4.089152753e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.41 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.412257709e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -3.015082478e-8   k1 = 4.681262989e-01 wk1 = 1.082750080e-7   k2 = -4.122919261e-02 wk2 = -2.617090033e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.319130474e+05 wvsat = 1.140986381e-1   ua = -1.249558358e-09 wua = 4.496676663e-16   ub = 2.609314994e-18 wub = -3.773118814e-25   uc = 1.264656591e-10 wuc = -1.730756901e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.260217473e-02 wu0 = -5.560639416e-10   a0 = 1.387952274e+00 wa0 = 8.952614623e-7   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 5.672929384e-01 wags = -1.315732378e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.204319435e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.695240176e-8   nfactor = {8.491646233e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.177733710e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.156851852e-06 wcit = 1.854659268e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 5.655476770e-03 wpdiblc2 = 3.181111576e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.523936430e-05 walpha0 = 1.079791528e-11   alpha1 = 0.0   beta0 = 1.779868928e+01 wbeta0 = -8.854143344e-9   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.535465922e-01 wkt1 = -6.788052919e-9   kt2 = -3.282950933e-02 wkt2 = -5.875560560e-9   at = 6.389441389e+05 wat = -9.653501488e-1   ute = -1.359755904e+00 wute = 2.974873465e-7   ua1 = 2.234265226e-09 wua1 = -4.499403383e-16   ub1 = -2.855474330e-18 wub1 = 2.309792652e-24   uc1 = -1.825682696e-10 wuc1 = 4.089152753e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.42 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.397854649e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.676677975e-09 wvth0 = -3.782482399e-08 pvth0 = 3.024553307e-14   k1 = 5.114861770e-01 lk1 = -1.708942876e-07 wk1 = 1.577451915e-07 pk1 = -1.949768342e-13   k2 = -6.374524485e-02 lk2 = 8.874251668e-08 wk2 = -3.691128402e-08 pk2 = 4.233107423e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.284401914e+05 lvsat = -3.804424325e-01 wvsat = 2.083404178e-01 pvsat = -3.714351263e-7   ua = -1.114226441e-09 lua = -5.333836831e-16 wua = 4.357639884e-16 pua = 5.479856564e-23   ub = 2.561792756e-18 lub = 1.872993957e-25 wub = -5.940949781e-25 pub = 8.544072189e-31   uc = 1.181571877e-10 luc = 3.274617835e-17 wuc = -2.062419557e-16 puc = 1.307182026e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.427590413e-02 lu0 = -6.596669665e-09 wu0 = -3.550558237e-09 pu0 = 1.180220037e-14   a0 = 9.194582417e-01 la0 = 1.846475528e-06 wa0 = 1.810750413e-06 pa0 = -3.608216603e-12   keta = 3.287786852e-01 lketa = -1.295815432e-06 wketa = -2.541197636e-07 pketa = 1.001562224e-12   a1 = 0.0   a2 = 0.38689047   ags = -1.055052769e+00 lags = 6.394151138e-06 wags = 1.042058260e-06 pags = -4.625633821e-12   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.218552076e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.609510935e-09 wvoff = 3.029973810e-08 pvoff = -5.260585673e-14   nfactor = {5.079280551e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.344915687e-06 wnfactor = 2.063678736e-06 pnfactor = -3.491775132e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.156851852e-06 wcit = 1.854659268e-11   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374771338e-01 letab = 2.659476276e-07 wetab = 2.819152378e-11 petab = -1.111112527e-16   dsub = 8.387771218e-01 ldsub = -1.098744270e-06 wdsub = -2.088748882e-07 pdsub = 8.232385968e-13   voffl = 0.0   minv = 0.0   pclm = 2.764451653e-01 lpclm = -3.012933301e-07 wpclm = -1.827948483e-07 ppclm = 7.204493357e-13   pdiblc1 = 0.39   pdiblc2 = 7.896089392e-03 lpdiblc2 = -8.830926525e-09 wpdiblc2 = -7.286476814e-09 ppdiblc2 = 4.125590612e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.940740981e-05 lalpha0 = 4.912703308e-10 walpha0 = 8.456315792e-11 palpha0 = -2.907309508e-16   alpha1 = 0.0   beta0 = 1.390340098e+01 lbeta0 = 1.535249980e-05 wbeta0 = 9.838079339e-07 pbeta0 = -3.912379045e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.716308015e-01 lkt1 = 7.127529399e-08 wkt1 = 4.084590106e-08 pkt1 = -1.877397028e-13   kt2 = -3.052087126e-02 lkt2 = -9.099035228e-09 wkt2 = -8.543494037e-09 pkt2 = 1.051512621e-14   at = 1.225365560e+06 lat = -2.311262746e+00 wat = -1.925572171e+00 pat = 3.784523057e-6   ute = -1.396537470e+00 lute = 1.449671886e-07 wute = 2.600426661e-07 pute = 1.475807188e-13   ua1 = 2.021873812e-09 lua1 = 8.370982786e-16 wua1 = -2.303128861e-16 pua1 = -8.656176774e-22   ub1 = -2.477214653e-18 lub1 = -1.490834865e-24 wub1 = 2.372080437e-24 pub1 = -2.454948495e-31   uc1 = -2.549182016e-10 luc1 = 2.851527868e-16 wuc1 = 6.463437125e-16 puc1 = -9.357766997e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.43 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.446122559e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.693571407e-09 wvth0 = -3.092953368e-08 pvth0 = 1.685970599e-14   k1 = 4.329315891e-01 lk1 = -1.839626604e-08 wk1 = 4.226025494e-08 pk1 = 2.921407320e-14   k2 = -1.759972644e-02 lk2 = -8.397782177e-10 wk2 = -7.368689256e-09 pk2 = -1.501996498e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3.635840048e+03 lvsat = 7.008676729e-02 wvsat = 1.224470827e-02 pvsat = 9.245474673e-9   ua = -1.319860560e-09 lua = -1.341861681e-16 wua = 9.718871926e-16 pua = -9.859774105e-22   ub = 2.653811067e-18 lub = 8.664248595e-27 wub = -4.494314421e-25 pub = 5.735718965e-31   uc = 1.593155388e-10 luc = -4.715452870e-17 wuc = -1.684383571e-16 puc = 5.733007682e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.251184299e-02 lu0 = -3.172097771e-09 wu0 = 7.245439540e-09 pu0 = -9.156070119e-15   a0 = 2.040146365e+00 la0 = -3.291163253e-07 wa0 = 3.113706904e-07 pa0 = -6.974707466e-13   keta = -3.984493389e-01 lketa = 1.159523311e-07 wketa = 2.535635698e-07 pketa = 1.599656908e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.905639409e+00 lags = 6.465594119e-07 wags = -1.112995875e-06 pags = -4.420272286e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.205618863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.098786294e-09 wvoff = 2.898231878e-09 pvoff = 5.886872986e-16   nfactor = {6.176100235e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.131990081e-06 wnfactor = 6.452011943e-07 pnfactor = -7.380846799e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.952296500e-06 lcit = 1.125069670e-11 wcit = 3.600450036e-11 pcit = -3.389103619e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 4.947097019e-04 leta0 = 1.027005569e-11 weta0 = 1.128828311e-10 peta0 = -2.191394400e-16   etab = -4.907591150e-04 letab = 1.597834523e-11 wetab = -5.931597606e-11 petab = 5.876705675e-17   dsub = -4.559497036e-01 ldsub = 1.414708916e-06 wdsub = 1.159841333e-06 pdsub = -1.833850204e-12   voffl = 0.0   minv = 0.0   pclm = 2.918847761e-01 lpclm = -3.312662465e-07 wpclm = -5.996426108e-08 ppclm = 4.819983167e-13   pdiblc1 = 0.39   pdiblc2 = -4.255699307e-03 lpdiblc2 = 1.475934088e-08 wpdiblc2 = 2.199550173e-08 ppdiblc2 = -1.558919883e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.729653474e-04 lalpha0 = -2.122039028e-10 walpha0 = -1.258335773e-10 palpha0 = 1.177122312e-16   alpha1 = 0.0   beta0 = 2.270680122e+01 lbeta0 = -1.737541090e-06 wbeta0 = -1.864867576e-06 pbeta0 = 1.617754722e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.114486799e-01 lkt1 = -4.555625866e-08 wkt1 = -9.329209122e-08 pkt1 = 7.266238159e-14   kt2 = -5.067780126e-02 lkt2 = 3.003161298e-08 wkt2 = 9.577423365e-11 pkt2 = -6.256285281e-15   at = -3.419971708e+03 lat = 7.417860599e-02 wat = 4.145175518e-02 pat = -3.406049137e-8   ute = -1.509239021e+00 lute = 3.637547087e-07 wute = 6.056143540e-07 pute = -5.232775988e-13   ua1 = 1.405029824e-09 lua1 = 2.034577513e-15 wua1 = 1.145349319e-15 pua1 = -3.536190716e-21   ub1 = -1.873415519e-18 lub1 = -2.662990123e-24 wub1 = -2.986940249e-25 pub1 = 4.939279614e-30   uc1 = -8.315996621e-11 luc1 = -4.828147551e-17 wuc1 = 1.867546314e-16 puc1 = -4.357641651e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.44 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.538000940e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.234208341e-08 wvth0 = -1.656290742e-08 pvth0 = 3.336400696e-15   k1 = 4.435474899e-01 lk1 = -2.838901348e-08 wk1 = 5.513085952e-10 pk1 = 6.847470439e-14   k2 = -3.244500138e-02 lk2 = 1.313407908e-08 wk2 = 1.785400918e-08 pk2 = -3.876209102e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -4.807333056e+03 lvsat = 7.118949366e-02 wvsat = 5.141020457e-02 pvsat = -2.762100700e-8   ua = -2.284638170e-09 lua = 7.739589958e-16 wua = 1.782127078e-15 pua = -1.748656215e-21   ub = 3.646722621e-18 lub = -9.259633970e-25 wub = -1.530933767e-24 pub = 1.591590035e-30   uc = 1.720669607e-10 luc = -5.915744217e-17 wuc = -2.299453706e-16 puc = 1.152266285e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.605785733e-02 lu0 = 2.903038922e-09 wu0 = 1.011221689e-08 pu0 = -1.185456764e-14   a0 = 6.880373489e-01 la0 = 9.436238914e-07 wa0 = 1.902904923e-06 pa0 = -2.195581920e-12   keta = -4.943804739e-01 lketa = 2.062523085e-07 wketa = 4.697288230e-07 pketa = -1.874797838e-13   a1 = 0.0   a2 = 0.38689047   ags = 3.535230247e+00 lags = -8.873744440e-07 wags = -1.075083339e-06 pags = -4.777142991e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.353868111e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.705348794e-08 wvoff = 4.490584349e-08 pvoff = -3.895307751e-14   nfactor = {1.256307174e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.307844534e-07 wnfactor = -3.426496079e-07 pnfactor = 1.917792803e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.877607945e-03 leta0 = -3.174052060e-09 weta0 = -9.065667441e-09 peta0 = 8.420629931e-15   etab = -8.320534746e-04 letab = 3.372387260e-10 wetab = 8.970158400e-11 petab = -8.150317253e-17   dsub = 1.088446920e+00 ldsub = -3.903162584e-08 wdsub = -1.484183114e-06 pdsub = 6.549700083e-13   voffl = 0.0   minv = 0.0   pclm = -3.392820136e-01 lpclm = 2.628510526e-07 wpclm = 7.506008881e-07 ppclm = -2.809866583e-13   pdiblc1 = 0.39   pdiblc2 = 7.992103178e-03 lpdiblc2 = 3.230484397e-09 wpdiblc2 = 2.191926845e-08 ppdiblc2 = -1.551744044e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.660419144e-05 lalpha0 = 1.969585332e-11 walpha0 = -1.035899462e-10 palpha0 = 9.677430126e-17   alpha1 = 0.0   beta0 = 1.890049540e+01 lbeta0 = 1.845334576e-06 wbeta0 = -2.039375194e-06 pbeta0 = 1.782018743e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.745073462e-01 lkt1 = 1.380086394e-08 wkt1 = 9.961360089e-09 pkt1 = -2.453009212e-14   kt2 = -2.516567694e-02 lkt2 = 6.017050355e-09 wkt2 = 2.327079337e-08 pkt2 = -2.807093080e-14   at = 8.885696405e+04 lat = -1.268167364e-02 wat = -2.130001612e-02 pat = 2.500775095e-8   ute = -3.035898097e-01 lute = -7.711228938e-07 wute = -1.258850794e-06 pute = 1.231743445e-12   ua1 = 7.721065106e-09 lua1 = -3.910706498e-15 wua1 = -8.733220368e-15 pua1 = 5.762506930e-21   ub1 = -1.012715536e-17 lub1 = 5.106255193e-24 wub1 = 1.333029865e-23 pub1 = -7.889691188e-30   uc1 = -2.658420719e-10 luc1 = 1.236771905e-16 wuc1 = 3.027550603e-16 puc1 = -1.527676202e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.45 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.994549725e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.248958127e-08 wvth0 = -1.559840670e-08 pvth0 = 2.910766530e-15   k1 = 2.274643583e-01 lk1 = 6.696847247e-08 wk1 = 2.456468187e-07 pk1 = -3.968594424e-14   k2 = 4.184259104e-02 lk2 = -1.964903545e-08 wk2 = -1.123255584e-07 pk2 = 1.868615213e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.566093962e+05 lvsat = -4.370896658e-05 wvsat = 4.142432870e-03 pvsat = -6.761739346e-9   ua = 6.776669596e-10 lua = -5.333062578e-16 wua = -3.755989206e-15 pua = 6.953145014e-22   ub = 4.506546096e-19 lub = 4.844614165e-25 wub = 3.642272974e-24 pub = -6.913460999e-31   uc = 2.540302271e-11 luc = 5.565353682e-18 wuc = 7.112025075e-17 puc = -1.763363014e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.119538843e-02 lu0 = -3.777153548e-09 wu0 = -2.778616260e-08 pu0 = 4.869987232e-15   a0 = 3.864396664e+00 la0 = -4.581034745e-07 wa0 = -5.480547988e-06 pa0 = 1.062735850e-12   keta = -1.646581149e-02 lketa = -4.651431973e-09 wketa = 6.185210931e-08 pketa = -7.483790017e-15   a1 = 0.0   a2 = 0.38689047   ags = 2.690890656e+00 lags = -5.147673825e-07 wags = -3.808594306e-06 pags = 7.285840908e-13   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.692572027e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.332391424e-09 wvoff = -7.393477531e-08 pvoff = 1.349128757e-14   nfactor = {2.418012080e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.812407838e-08 wnfactor = 4.582258075e-07 pnfactor = -1.616470406e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 9.711223037e-06 lcit = -2.079062726e-12 wcit = -1.419185272e-11 pcit = 6.262864603e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.716055463e-02 leta0 = 6.110089083e-09 weta0 = 3.283002897e-08 peta0 = -1.006794089e-14   etab = 2.354465226e-02 letab = -1.042020151e-08 wetab = -2.855787988e-08 petab = 1.256067453e-14   dsub = 1.643321849e+00 ldsub = -2.838979321e-07 wdsub = -2.417916470e-07 pdsub = 1.067026538e-13   voffl = 0.0   minv = 0.0   pclm = 3.603742536e-01 lpclm = -4.590725805e-08 wpclm = -3.566197723e-07 ppclm = 2.076298192e-13   pdiblc1 = 0.39   pdiblc2 = 9.441160004e-03 lpdiblc2 = 2.591015619e-09 wpdiblc2 = -9.804781148e-09 ppdiblc2 = -1.517617351e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.971883945e-03 lalpha0 = 9.016286680e-10 walpha0 = 1.890465649e-09 palpha0 = -7.832024328e-16   alpha1 = 0.0   beta0 = 1.692195698e+01 lbeta0 = 2.718463582e-06 wbeta0 = 5.055179170e-06 pbeta0 = -1.348808098e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.221873536e-01 lkt1 = -9.287948805e-09 wkt1 = -7.991213414e-08 pkt1 = 1.513108088e-14   kt2 = -1.171197684e-02 lkt2 = 7.993249841e-11 wkt2 = -5.442567208e-08 pkt2 = 6.216519405e-15   at = 5.991169541e+04 lat = 9.187341105e-05 wat = 7.165691963e-02 pat = -1.601414479e-8   ute = -1.693087989e+00 lute = -1.579373473e-07 wute = 7.986007015e-07 pute = 3.237901000e-13   ua1 = -9.634638931e-10 lua1 = -7.822385072e-17 wua1 = 4.440625470e-15 pua1 = -5.111123803e-23   ub1 = 1.632196801e-18 lub1 = -8.314691739e-26 wub1 = -5.411955712e-24 pub1 = 3.812656610e-31   uc1 = 8.373378192e-11 luc1 = -3.059063373e-17 wuc1 = -1.827358888e-16 puc1 = 6.147953564e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.46 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.717341158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.718658138e-08 wvth0 = 2.375189569e-07 pvth0 = -4.551058513e-14   k1 = 4.593817134e-01 lk1 = 2.260268245e-08 wk1 = -1.392992291e-07 pk1 = 3.395423471e-14   k2 = -6.792606655e-02 lk2 = 1.349708746e-09 wk2 = 3.548579196e-08 pk2 = -9.590159181e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.667456932e+05 lvsat = -1.982782579e-03 wvsat = -3.786474290e-02 pvsat = 1.274233378e-9   ua = -2.036253991e-09 lua = -1.413317991e-17 wua = -4.963000267e-17 pua = -1.371201421e-23   ub = 3.290750186e-18 lub = -5.884886720e-26 wub = 8.028519546e-25 pub = -1.481648589e-31   uc = 6.399617735e-11 luc = -1.817516802e-18 wuc = -5.245744757e-18 puc = -3.024815199e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.908352713e-02 lu0 = -1.460154483e-09 wu0 = 6.744966381e-09 pu0 = -1.735817742e-15   a0 = 4.016508677e+00 la0 = -4.872025025e-07 wa0 = 2.043859943e-07 pa0 = -2.479202111e-14   keta = 9.812353272e-02 lketa = -2.657237352e-08 wketa = 1.013667880e-08 pketa = 2.409371839e-15   a1 = 0.0   a2 = 0.38689047   ags = -2.078344509e+00 lags = 3.975873045e-07 wags = 3.021027986e-07 pags = -5.779226537e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.298462295e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.878301996e-09 wvoff = -3.780750763e-08 pvoff = 6.580141261e-15   nfactor = {2.747963881e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.499570108e-08 wnfactor = -3.234745567e-06 pnfactor = 5.448183834e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.182579656e-05 lcit = 2.040969123e-12 wcit = 5.068518827e-11 pcit = -6.148113337e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.109419257e-01 leta0 = 2.405046536e-08 weta0 = -1.676767560e-08 peta0 = -5.799000099e-16   etab = -6.988481150e-02 letab = 7.452854902e-09 wetab = 1.346421485e-07 petab = -1.865949090e-14   dsub = -1.385898727e-01 ldsub = 5.698178031e-08 wdsub = 8.412711567e-07 pdsub = -1.004872605e-13   voffl = 0.0   minv = 0.0   pclm = 3.160198970e-02 lpclm = 1.698687603e-08 wpclm = 1.784641104e-06 ppclm = -2.019933864e-13   pdiblc1 = -6.555542783e-01 lpdiblc1 = 2.000145334e-07 wpdiblc1 = -1.909803905e-08 ppdiblc1 = 3.653454869e-15   pdiblc2 = 4.593493264e-02 lpdiblc2 = -4.390243087e-09 wpdiblc2 = -6.190281930e-08 ppdiblc2 = 8.448737348e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 6.392563525e-03 lalpha0 = -6.984901330e-10 walpha0 = -5.555418537e-09 palpha0 = 6.411952120e-16   alpha1 = 0.0   beta0 = 3.478162342e+01 lbeta0 = -6.980906095e-07 wbeta0 = -3.483527987e-06 pbeta0 = 2.846465809e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.194027583e-01 lkt1 = -9.820641879e-09 wkt1 = 8.761251409e-09 pkt1 = -1.832137774e-15   kt2 = 9.064114085e-03 lkt2 = -3.894533695e-09 wkt2 = -6.622290363e-08 pkt2 = 8.473329801e-15   at = 5.063776336e+04 lat = 1.865976613e-03 wat = -5.603373945e-02 pat = 8.413078291e-9   ute = -3.972679210e+00 lute = 2.781484532e-07 wute = 7.038146833e-06 pute = -8.698350749e-13   ua1 = -4.163191824e-09 lua1 = 5.338841025e-16 wua1 = 1.277862669e-14 pua1 = -1.646170872e-21   ub1 = 3.325414154e-18 lub1 = -4.070593968e-25 wub1 = -1.070702586e-23 pub1 = 1.394212580e-30   uc1 = -1.622616570e-10 luc1 = 1.646829373e-17 wuc1 = 2.717790613e-16 puc1 = -2.546917431e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.47 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.819687682e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.842804472e-08 wvth0 = -5.000948379e-07 pvth0 = 4.396196818e-14   k1 = 6.380761762e-01 lk1 = 9.270441155e-10 wk1 = 5.685746075e-07 pk1 = -5.191086167e-14   k2 = -1.477594291e-01 lk2 = 1.103349562e-08 wk2 = -1.231906748e-07 pk2 = 9.657296236e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.019119850e+05 lvsat = -6.248453771e-03 wvsat = -1.183693744e-01 pvsat = 1.103944518e-8   ua = -2.077494297e-09 lua = -9.130730730e-18 wua = 3.709450189e-16 pua = -6.472776433e-23   ub = 4.150779493e-18 lub = -1.631704222e-25 wub = -2.708217801e-24 pub = 2.777279025e-31   uc = 1.135639425e-10 luc = -7.830086714e-18 wuc = -1.220374679e-16 puc = 1.114202082e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.109570636e-02 lu0 = -1.704231824e-09 wu0 = -2.325418033e-08 pu0 = 1.903078753e-15   a0 = 0.0   keta = 4.637224546e-02 lketa = -2.029494237e-08 wketa = 1.212983659e-07 pketa = -1.107454081e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.053216521e+00 lags = 1.772895167e-08 wags = -7.049065300e-07 pags = 6.435796619e-14   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.450772724e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.725827491e-09 wvoff = 6.646968618e-08 pvoff = -6.068682348e-15   nfactor = {4.091164824e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.833697347e-07 wnfactor = 1.168797299e-06 pnfactor = 1.066863375e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.021666667e-05 lcit = 1.845781667e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.122598964e-01 leta0 = -3.023915659e-09 weta0 = -8.712730200e-08 peta0 = 7.954722672e-15   etab = -3.413909109e-02 letab = 3.116899017e-09 wetab = -7.757994297e-08 petab = 7.083048793e-15   dsub = 5.477609584e-01 ldsub = -2.627257550e-08 wdsub = 5.196435957e-08 pdsub = -4.744346029e-15   voffl = 0.0   minv = 0.0   pclm = 1.826961459e-01 lpclm = -1.340845122e-09 wpclm = 4.827859830e-07 ppclm = -4.407836025e-14   pdiblc1 = 9.731933160e-01 lpdiblc1 = 2.447450247e-09 wpdiblc1 = 4.456209111e-08 ppdiblc1 = -4.068518918e-15   pdiblc2 = 2.163491443e-02 lpdiblc2 = -1.442650878e-09 wpdiblc2 = 3.133084556e-08 ppdiblc2 = -2.860506199e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.546768328e-03 lalpha0 = -1.106951756e-10 walpha0 = -1.089235218e-09 palpha0 = 9.944717544e-17   alpha1 = 0.0   beta0 = 3.226222131e+01 lbeta0 = -3.924871334e-07 wbeta0 = -4.596845462e-06 pbeta0 = 4.196919907e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.317769488e-01 lkt1 = -2.044965258e-08 wkt1 = -2.564659928e-08 pkt1 = 2.341534515e-15   kt2 = -5.771372187e-02 lkt2 = 4.205617807e-09 wkt2 = 1.468305304e-08 pkt2 = -1.340562743e-15   at = 1.909806949e+03 lat = 7.776677726e-03 wat = 5.387285651e-02 pat = -4.918591799e-9   ute = -1.728970497e+00 lute = 5.986586382e-09 wute = -5.369288037e-07 pute = 4.902159978e-14   ua1 = 4.973649069e-10 lua1 = -3.144142900e-17 wua1 = -3.204115137e-15 pua1 = 2.925357120e-22   ub1 = 1.190106824e-19 lub1 = -1.812265580e-26 wub1 = 3.181678112e-24 pub1 = -2.904872117e-31   uc1 = 1.218817138e-11 luc1 = -4.692470447e-18 wuc1 = 2.499208607e-16 puc1 = -2.281777458e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.48 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.49 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.50 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.170316381e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.387112143e-8   k1 = 6.063790645e-01 lk1 = -2.881841689e-7   k2 = -8.594952435e-02 lk2 = 1.142071145e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.537690438e+05 lvsat = -6.038822173e-1   ua = -8.520891125e-10 lua = -5.004191656e-16   ub = 2.204410149e-18 lub = 7.012749237e-25   uc = -5.909317978e-12 luc = 1.113807635e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214003729e-02 lu0 = 5.030387991e-10   a0 = 2.008729703e+00 la0 = -3.240761624e-7   keta = 1.759108995e-01 lketa = -6.933176282e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.281942499e-01 lags = 3.611563944e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.036281567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.603596488e-8   nfactor = {1.749350581e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.555897014e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 7.131267544e-01 ldsub = -6.035184771e-7   voffl = 0.0   minv = 0.0   pclm = 1.664834555e-01 lpclm = 1.320987568e-7   pdiblc1 = 0.39   pdiblc2 = 3.512850715e-03 lpdiblc2 = 1.598689531e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.853776267e-05 lalpha0 = 3.163787912e-10 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.449521854e+01 lbeta0 = 1.299897675e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470596215e-01 lkt1 = -4.166103278e-8   kt2 = -3.566027875e-02 lkt2 = -2.773576563e-9   at = 6.702214770e+04 lat = -3.465249173e-2   ute = -1.240106715e+00 lute = 2.337455558e-7   ua1 = 1.883327245e-09 lua1 = 3.163790093e-16   ub1 = -1.050270605e-18 lub1 = -1.638514265e-24   uc1 = 1.338950523e-10 luc1 = -2.777712061e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.51 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.260063464e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.448520205e-9   k1 = 4.583535850e-01 lk1 = -8.223055605e-10   k2 = -2.203242067e-02 lk2 = -9.875158843e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.730062600e+03 lvsat = 7.564845687e-2   ua = -7.352140101e-10 lua = -7.273088020e-16   ub = 2.383451972e-18 lub = 3.537010318e-25   uc = 5.799009160e-11 luc = -1.266716032e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.687039536e-02 lu0 = -8.680005323e-9   a0 = 2.227453906e+00 la0 = -7.486854573e-7   keta = -2.459161360e-01 lketa = 1.255751958e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.236107797e+00 lags = 3.806543807e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.188184317e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.452915869e-9   nfactor = {1.005735986e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.879893114e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.470650000e-05 lcit = -9.136728450e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.626152760e-04 leta0 = -1.215550353e-10   etab = -5.264411170e-04 letab = 5.133014043e-11   dsub = 2.417621702e-01 ldsub = 3.115415901e-7   voffl = 0.0   minv = 0.0   pclm = 2.558127930e-01 lpclm = -4.131628605e-8   pdiblc1 = 0.39   pdiblc2 = 8.975871500e-03 lpdiblc2 = 5.381533057e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.972691479e-04 lalpha0 = -1.413931643e-10   alpha1 = 0.0   beta0 = 2.158497514e+01 lbeta0 = -7.643677381e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675692870e-01 lkt1 = -1.845619147e-9   kt2 = -5.062018750e-02 lkt2 = 2.626809429e-8   at = 2.151566470e+04 lat = 5.368924372e-2   ute = -1.144926840e+00 lute = 4.897286449e-8   ua1 = 2.094023910e-09 lua1 = -9.264642648e-17   ub1 = -2.053097310e-18 lub1 = 3.082732179e-25   uc1 = 2.918378297e-11 luc1 = -7.449521901e-17 wuc1 = -6.162975822e-33 puc1 = -1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.52 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.438365440e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.033504477e-8   k1 = 4.438791340e-01 lk1 = 1.280249517e-8   k2 = -2.170477869e-02 lk2 = -1.018356824e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.611888860e+04 lvsat = 5.457385496e-2   ua = -1.212585306e-09 lua = -2.779592013e-16   ub = 2.725777112e-18 lub = 3.147037747e-26   uc = 3.374147540e-11 luc = 1.015806211e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214094266e-02 lu0 = -4.228171494e-9   a0 = 1.832745096e+00 la0 = -3.771460549e-7   keta = -2.118113260e-01 lketa = 9.347233816e-8   a1 = 0.0   a2 = 0.38689047   ags = 2.888505226e+00 lags = -1.174747319e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.083733401e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.379048837e-9   nfactor = {1.050183549e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.461508205e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.575917150e-03 leta0 = 1.891445537e-9   etab = -7.780927660e-04 letab = 2.882098376e-10   dsub = 1.956246419e-01 ldsub = 3.549708455e-7   voffl = 0.0   minv = 0.0   pclm = 1.122479820e-01 lpclm = 9.382127054e-8   pdiblc1 = 0.39   pdiblc2 = 2.117781524e-02 lpdiblc2 = -6.104156585e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.571117306e-05 lalpha0 = 7.791121185e-11   alpha1 = 0.0   beta0 = 1.767369287e+01 lbeta0 = 2.917322269e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.685150100e-01 lkt1 = -9.554100870e-10   kt2 = -1.116694420e-02 lkt2 = -1.086924362e-8   at = 7.604376820e+04 lat = 2.361939893e-3   ute = -1.060861620e+00 lute = -3.015772709e-8   ua1 = 2.467526220e-09 lua1 = -4.442241509e-16   ub1 = -2.108207100e-18 lub1 = 3.601480632e-25   uc1 = -8.371733260e-11 luc1 = 3.177860108e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.53 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.900716256e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.073858628e-8   k1 = 3.752351760e-01 lk1 = 4.309507383e-8   k2 = -2.572775116e-02 lk2 = -8.408230486e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.591013100e+05 lvsat = -4.111287603e-3   ua = -1.581778528e-09 lua = -1.150342324e-16   ub = 2.641693184e-18 lub = 6.857661490e-26   uc = 6.818598102e-11 luc = -5.042298220e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.448039904e-02 lu0 = -8.475735971e-10   a0 = 5.675289840e-01 la0 = 1.811938154e-7   keta = 2.074182187e-02 lketa = -9.153365992e-9   a1 = 0.0   a2 = 0.38689047   ags = 3.998001480e-01 lags = -7.648176831e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.314017785e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.783401020e-9   nfactor = {2.693661497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.911599775e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.174000000e-06 lcit = 1.688413800e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.588613096e-03 leta0 = 5.363834004e-11   etab = 6.365430149e-03 letab = -2.864226825e-09 wetab = 1.344168495e-24 petab = -1.232595164e-32   dsub = 1.497870141e+00 ldsub = -2.197100933e-7   voffl = 0.0   minv = 0.0   pclm = 1.458467640e-01 lpclm = 7.899412805e-8   pdiblc1 = 0.39   pdiblc2 = 3.543015120e-03 lpdiblc2 = 1.678080708e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.346591437e-04 lalpha0 = 4.304869513e-10 palpha0 = 4.930380658e-32   alpha1 = 0.0   beta0 = 1.996294063e+01 lbeta0 = 1.907077232e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702591400e-01 lkt1 = -1.857255180e-10   kt2 = -4.445217720e-02 lkt2 = 3.819529698e-9   at = 1.030174912e+05 lat = -9.541564067e-3   ute = -1.212683320e+00 lute = 3.684118912e-8   ua1 = 1.707830040e-09 lua1 = -1.089702267e-16   ub1 = -1.623408644e-18 lub1 = 1.462065046e-25   uc1 = -2.619246032e-11 luc1 = 6.392874939e-18 wuc1 = 6.162975822e-33   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.54 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.146155529e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.456383956e-8   k1 = 3.755851429e-01 lk1 = 4.302812517e-8   k2 = -4.657930326e-02 lk2 = -4.419328570e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.439678529e+05 lvsat = -1.216257252e-3   ua = -2.066109318e-09 lua = -2.238175224e-17   ub = 3.773712230e-18 lub = -1.479786286e-25   uc = 6.084055744e-11 luc = -3.637118691e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.314101586e-02 lu0 = -2.504349593e-9   a0 = 4.139458714e+00 la0 = -5.021163420e-7   keta = 1.042213333e-01 lketa = -2.512299653e-08 wketa = -2.646977960e-23 pketa = -6.310887242e-30   a1 = 0.0   a2 = 0.38689047   ags = -1.896612143e+00 lags = 3.628219029e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.525896395e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.836638845e-9   nfactor = {8.020766929e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.827441752e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.866428571e-05 lcit = -1.657477857e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.210286556e-01 leta0 = 2.370162185e-08 weta0 = 2.316105715e-23 peta0 = -5.127595884e-30   etab = 1.111025482e-02 letab = -3.771911785e-9   dsub = 3.674835515e-01 ldsub = -3.467138701e-9   voffl = 0.0   minv = 0.0   pclm = 1.105167186e+00 lpclm = -1.045238686e-7   pdiblc1 = -6.670428571e-01 lpdiblc1 = 2.022122986e-7   pdiblc2 = 8.696794286e-03 lpdiblc2 = 6.921627531e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.050656864e-03 lalpha0 = -3.127740010e-10   alpha1 = 0.0   beta0 = 3.268607917e+01 lbeta0 = -5.268591715e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.141323571e-01 lkt1 = -1.092277908e-8   kt2 = -3.077280571e-02 lkt2 = 1.202665933e-9   at = 1.693021714e+04 lat = 6.926931461e-3   ute = 2.611745714e-01 lute = -2.451078255e-7   ua1 = 3.523893743e-09 lua1 = -4.563832130e-16   ub1 = -3.115483286e-18 lub1 = 4.316403836e-25 wub1 = 7.346839693e-40   uc1 = 1.229221143e-12 luc1 = 1.147107275e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.55 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.65e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.005206618e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.646412928e-08 wvth0 = -1.984645783e-07 pvth0 = 2.407375335e-14   k1 = 1.048218798e+00 lk1 = -3.856233722e-08 wk1 = -1.132259802e-07 pk1 = 1.373431140e-14   k2 = -2.361228856e-01 lk2 = 1.857230797e-08 wk2 = 2.370031721e-08 pk2 = -2.874848477e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 7.646281157e+04 lvsat = 6.972104257e-03 wvsat = 9.017105901e-02 pvsat = -1.093774946e-8   ua = -4.222622995e-10 lua = -2.217803956e-16 wua = -2.380629893e-15 pua = 2.887704060e-22   ub = 1.949692343e-18 lub = 7.327498371e-26 wub = 9.507594229e-25 pub = -1.153271180e-31   uc = -4.582367333e-11 luc = 9.301252501e-18 wuc = 1.429205352e-16 puc = -1.733626092e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.133133105e-02 lu0 = -2.284834827e-09 wu0 = -2.364587103e-08 pu0 = 2.868244156e-15   a0 = 0.0   keta = 9.531613622e-01 lketa = -1.280994220e-07 wketa = -1.386102522e-06 pketa = 1.681342359e-13   a1 = 0.0   a2 = 0.38689047   ags = 6.215905339e-01 lags = 5.736391823e-08 wags = 1.260692891e-08 pags = -1.529220476e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.499221232e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.964306912e-08 wvoff = 2.407585240e-07 pvoff = -2.920400897e-14   nfactor = {-2.315266125e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.608778591e-07 wnfactor = 5.085589421e-06 pnfactor = -6.168819968e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.021666667e-05 lcit = 1.845781667e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -8.766673793e-02 leta0 = 1.965482123e-08 weta0 = 2.452207386e-07 peta0 = -2.974527560e-14   etab = -1.361934351e-01 letab = 1.409602581e-08 wetab = 9.207009586e-08 petab = -1.116810263e-14   dsub = 5.790205365e-01 ldsub = -2.912657498e-8   voffl = 0.0   minv = 0.0   pclm = 1.242638577e+00 lpclm = -1.211991484e-07 wpclm = -1.279209318e-06 ppclm = 1.551680902e-13   pdiblc1 = 7.629136521e-01 lpdiblc1 = 2.875857400e-08 wpdiblc1 = 3.941204905e-07 ppdiblc1 = -4.780681549e-14   pdiblc2 = 4.856372255e-02 lpdiblc2 = -4.143695646e-09 wpdiblc2 = -1.343425862e-08 ppdiblc2 = 1.629575570e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.874307615e-04 lalpha0 = 3.453532524e-11 walpha0 = 1.170459585e-09 palpha0 = -1.419767477e-16   alpha1 = 0.0   beta0 = 2.439057131e+01 lbeta0 = 4.793859325e-07 wbeta0 = 8.488591924e-06 pbeta0 = -1.029666200e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 1.498430755e-01 lkt1 = -5.507299906e-08 wkt1 = -4.937976466e-07 pkt1 = 5.989765454e-14   kt2 = -3.122450640e-02 lkt2 = 1.257457227e-09 wkt2 = -2.935129429e-08 pkt2 = 3.560311998e-15   at = -2.870865609e+04 lat = 1.246292678e-02 wat = 1.047714585e-01 pat = -1.270877792e-8   ute = -2.008831474e+00 lute = 3.024390784e-08 wute = -7.170190816e-08 pute = 8.697441460e-15   ua1 = -2.681328401e-09 lua1 = 2.963102330e-16 wua1 = 2.079985683e-15 pua1 = -2.523022634e-22   ub1 = 4.186370853e-18 lub1 = -4.540745234e-25 wub1 = -3.579698066e-24 pub1 = 4.342173755e-31   uc1 = 2.862408008e-10 luc1 = -3.342479734e-17 wuc1 = -2.056505278e-16 puc1 = 2.494540902e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.56 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.57 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.58 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.170316381e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.387112143e-8   k1 = 6.063790645e-01 lk1 = -2.881841689e-7   k2 = -8.594952435e-02 lk2 = 1.142071145e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.537690438e+05 lvsat = -6.038822173e-1   ua = -8.520891125e-10 lua = -5.004191656e-16   ub = 2.204410149e-18 lub = 7.012749237e-25   uc = -5.909317978e-12 luc = 1.113807635e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214003729e-02 lu0 = 5.030387991e-10   a0 = 2.008729703e+00 la0 = -3.240761624e-7   keta = 1.759108995e-01 lketa = -6.933176282e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.281942499e-01 lags = 3.611563944e-06 pags = 1.615587134e-27   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.036281567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.603596488e-8   nfactor = {1.749350581e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.555897014e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 7.131267544e-01 ldsub = -6.035184771e-7   voffl = 0.0   minv = 0.0   pclm = 1.664834555e-01 lpclm = 1.320987568e-7   pdiblc1 = 0.39   pdiblc2 = 3.512850715e-03 lpdiblc2 = 1.598689531e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.853776267e-05 lalpha0 = 3.163787912e-10 palpha0 = 9.860761315e-32   alpha1 = 0.0   beta0 = 1.449521854e+01 lbeta0 = 1.299897675e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470596215e-01 lkt1 = -4.166103278e-8   kt2 = -3.566027875e-02 lkt2 = -2.773576563e-9   at = 6.702214770e+04 lat = -3.465249173e-2   ute = -1.240106715e+00 lute = 2.337455558e-7   ua1 = 1.883327245e-09 lua1 = 3.163790093e-16   ub1 = -1.050270605e-18 lub1 = -1.638514265e-24   uc1 = 1.338950523e-10 luc1 = -2.777712061e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.59 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.260063464e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.448520205e-9   k1 = 4.583535850e-01 lk1 = -8.223055605e-10   k2 = -2.203242067e-02 lk2 = -9.875158843e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.730062600e+03 lvsat = 7.564845687e-2   ua = -7.352140101e-10 lua = -7.273088020e-16   ub = 2.383451972e-18 lub = 3.537010318e-25   uc = 5.799009160e-11 luc = -1.266716032e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.687039536e-02 lu0 = -8.680005323e-9   a0 = 2.227453906e+00 la0 = -7.486854573e-7   keta = -2.459161360e-01 lketa = 1.255751958e-07 wketa = -2.117582368e-22   a1 = 0.0   a2 = 0.38689047   ags = 1.236107797e+00 lags = 3.806543807e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.188184317e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.452915869e-9   nfactor = {1.005735986e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.879893114e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.470650000e-05 lcit = -9.136728450e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.626152760e-04 leta0 = -1.215550353e-10   etab = -5.264411170e-04 letab = 5.133014043e-11   dsub = 2.417621702e-01 ldsub = 3.115415901e-7   voffl = 0.0   minv = 0.0   pclm = 2.558127930e-01 lpclm = -4.131628605e-8   pdiblc1 = 0.39   pdiblc2 = 8.975871500e-03 lpdiblc2 = 5.381533057e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.972691479e-04 lalpha0 = -1.413931643e-10   alpha1 = 0.0   beta0 = 2.158497514e+01 lbeta0 = -7.643677381e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675692870e-01 lkt1 = -1.845619147e-9   kt2 = -5.062018750e-02 lkt2 = 2.626809429e-8   at = 2.151566470e+04 lat = 5.368924372e-2   ute = -1.144926840e+00 lute = 4.897286449e-8   ua1 = 2.094023910e-09 lua1 = -9.264642648e-17   ub1 = -2.053097310e-18 lub1 = 3.082732179e-25   uc1 = 2.918378297e-11 luc1 = -7.449521901e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.60 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.438365440e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.033504477e-8   k1 = 4.438791340e-01 lk1 = 1.280249517e-8   k2 = -2.170477869e-02 lk2 = -1.018356824e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.611888860e+04 lvsat = 5.457385496e-2   ua = -1.212585306e-09 lua = -2.779592013e-16   ub = 2.725777112e-18 lub = 3.147037747e-26   uc = 3.374147540e-11 luc = 1.015806211e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214094266e-02 lu0 = -4.228171494e-9   a0 = 1.832745096e+00 la0 = -3.771460549e-7   keta = -2.118113260e-01 lketa = 9.347233816e-8   a1 = 0.0   a2 = 0.38689047   ags = 2.888505226e+00 lags = -1.174747319e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.083733401e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.379048837e-9   nfactor = {1.050183549e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.461508205e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.575917150e-03 leta0 = 1.891445537e-09 weta0 = 8.271806126e-25 peta0 = -7.888609052e-31   etab = -7.780927660e-04 letab = 2.882098376e-10   dsub = 1.956246419e-01 ldsub = 3.549708455e-7   voffl = 0.0   minv = 0.0   pclm = 1.122479820e-01 lpclm = 9.382127054e-8   pdiblc1 = 0.39   pdiblc2 = 2.117781524e-02 lpdiblc2 = -6.104156585e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.571117306e-05 lalpha0 = 7.791121185e-11 palpha0 = 2.465190329e-32   alpha1 = 0.0   beta0 = 1.767369287e+01 lbeta0 = 2.917322269e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.685150100e-01 lkt1 = -9.554100870e-10   kt2 = -1.116694420e-02 lkt2 = -1.086924362e-8   at = 7.604376820e+04 lat = 2.361939893e-3   ute = -1.060861620e+00 lute = -3.015772709e-8   ua1 = 2.467526220e-09 lua1 = -4.442241509e-16   ub1 = -2.108207100e-18 lub1 = 3.601480632e-25   uc1 = -8.371733260e-11 luc1 = 3.177860108e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.61 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.900716256e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.073858628e-8   k1 = 3.752351760e-01 lk1 = 4.309507383e-8   k2 = -2.572775116e-02 lk2 = -8.408230486e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.591013100e+05 lvsat = -4.111287603e-3   ua = -1.581778528e-09 lua = -1.150342324e-16   ub = 2.641693184e-18 lub = 6.857661490e-26   uc = 6.818598102e-11 luc = -5.042298220e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.448039904e-02 lu0 = -8.475735971e-10   a0 = 5.675289840e-01 la0 = 1.811938154e-7   keta = 2.074182187e-02 lketa = -9.153365992e-9   a1 = 0.0   a2 = 0.38689047   ags = 3.998001480e-01 lags = -7.648176831e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.314017785e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.783401020e-9   nfactor = {2.693661497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.911599775e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.174000000e-06 lcit = 1.688413800e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.588613096e-03 leta0 = 5.363834004e-11   etab = 6.365430149e-03 letab = -2.864226825e-09 wetab = 1.447566072e-24 petab = -3.451266460e-31   dsub = 1.497870141e+00 ldsub = -2.197100933e-7   voffl = 0.0   minv = 0.0   pclm = 1.458467640e-01 lpclm = 7.899412805e-8   pdiblc1 = 0.39   pdiblc2 = 3.543015120e-03 lpdiblc2 = 1.678080708e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.346591437e-04 lalpha0 = 4.304869513e-10 walpha0 = 4.135903063e-25   alpha1 = 0.0   beta0 = 1.996294063e+01 lbeta0 = 1.907077232e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702591400e-01 lkt1 = -1.857255180e-10   kt2 = -4.445217720e-02 lkt2 = 3.819529698e-9   at = 1.030174912e+05 lat = -9.541564067e-3   ute = -1.212683320e+00 lute = 3.684118912e-8   ua1 = 1.707830040e-09 lua1 = -1.089702267e-16   ub1 = -1.623408644e-18 lub1 = 1.462065046e-25   uc1 = -2.619246032e-11 luc1 = 6.392874939e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.62 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.146155529e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.456383956e-8   k1 = 3.755851429e-01 lk1 = 4.302812517e-8   k2 = -4.657930326e-02 lk2 = -4.419328570e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.439678529e+05 lvsat = -1.216257252e-3   ua = -2.066109318e-09 lua = -2.238175224e-17   ub = 3.773712230e-18 lub = -1.479786286e-25   uc = 6.084055744e-11 luc = -3.637118691e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.314101586e-02 lu0 = -2.504349593e-9   a0 = 4.139458714e+00 la0 = -5.021163420e-7   keta = 1.042213333e-01 lketa = -2.512299653e-08 wketa = 5.293955920e-23 pketa = -1.262177448e-29   a1 = 0.0   a2 = 0.38689047   ags = -1.896612143e+00 lags = 3.628219029e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.525896395e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.836638845e-9   nfactor = {8.020766929e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.827441752e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.866428571e-05 lcit = -1.657477857e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.210286556e-01 leta0 = 2.370162185e-08 weta0 = -6.617444900e-24 peta0 = 1.577721810e-30   etab = 1.111025482e-02 letab = -3.771911785e-9   dsub = 3.674835515e-01 ldsub = -3.467138701e-9   voffl = 0.0   minv = 0.0   pclm = 1.105167186e+00 lpclm = -1.045238686e-7   pdiblc1 = -6.670428571e-01 lpdiblc1 = 2.022122986e-07 ppdiblc1 = -1.009741959e-28   pdiblc2 = 8.696794286e-03 lpdiblc2 = 6.921627531e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.050656864e-03 lalpha0 = -3.127740010e-10   alpha1 = 0.0   beta0 = 3.268607917e+01 lbeta0 = -5.268591715e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.141323571e-01 lkt1 = -1.092277908e-8   kt2 = -3.077280571e-02 lkt2 = 1.202665933e-9   at = 1.693021714e+04 lat = 6.926931461e-3   ute = 2.611745714e-01 lute = -2.451078255e-7   ua1 = 3.523893743e-09 lua1 = -4.563832130e-16   ub1 = -3.115483286e-18 lub1 = 4.316403836e-25 wub1 = 1.469367939e-39 pub1 = -1.751623080e-46   uc1 = 1.229221143e-12 luc1 = 1.147107275e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.63 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-2.048011671e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.684128427e-07 wvth0 = 2.179072129e-06 pvth0 = -2.643214493e-13   k1 = 1.836162705e+00 lk1 = -1.341399331e-07 wk1 = -9.109009940e-07 pk1 = 1.104922906e-13   k2 = -5.377895772e-01 lk2 = 5.516447766e-08 wk2 = 3.290925925e-07 pk2 = -3.991893146e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.470174024e+05 lvsat = -1.371616761e-02 wvsat = -8.248988100e-02 pvsat = 1.000602257e-8   ua = -5.529489163e-09 lua = 3.977262230e-16 wua = 2.789671222e-15 pua = -3.383871193e-22   ub = 5.163859183e-18 lub = -3.166034540e-25 wub = -2.303102378e-24 pub = 2.793663184e-31   uc = 1.753861359e-11 luc = 1.615407098e-18 wuc = 7.877572405e-17 puc = -9.555495327e-24   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -2.793980063e-02 lu0 = 4.904753447e-09 wu0 = 3.635725913e-08 pu0 = -4.410135533e-15   a0 = 0.0   keta = -2.163891257e+00 lketa = 2.499990606e-07 wketa = 1.769445697e-06 pketa = -2.146337630e-13   a1 = 0.0   a2 = 0.38689047   ags = 5.902701670e-01 lags = 6.116307875e-08 wags = 4.431410241e-08 pags = -5.375300622e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {4.794227903e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.882646890e-08 wvoff = -4.975937992e-07 pvoff = 6.035812785e-14   nfactor = {1.253741917e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.140752867e-06 wnfactor = -9.950526538e-06 pnfactor = 1.206998869e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.021666667e-05 lcit = 1.845781667e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.509314225e-01 leta0 = 2.732882747e-08 weta0 = 3.092667420e-07 peta0 = -3.751405581e-14   etab = 1.105695349e-01 letab = -1.583632246e-08 wetab = -1.577403969e-07 petab = 1.913391014e-14   dsub = 5.796492536e-01 ldsub = -2.920283837e-08 wdsub = -6.364818116e-10 pdsub = 7.720524375e-17   voffl = 0.0   minv = 0.0   pclm = -2.680169996e-02 lpclm = 3.278395720e-08 wpclm = 5.908546988e-09 ppclm = -7.167067496e-16   pdiblc1 = 1.963163288e+00 lpdiblc1 = -1.168317069e-07 wpdiblc1 = -8.209522289e-07 ppdiblc1 = 9.958150536e-14   pdiblc2 = 2.170879397e-01 lpdiblc2 = -2.458568318e-08 wpdiblc2 = -1.840397498e-07 ppdiblc2 = 2.232402165e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.544942717e-03 lalpha0 = 2.446722282e-10 walpha0 = 2.924227876e-09 palpha0 = -3.547088414e-16   alpha1 = 0.0   beta0 = -6.913597331e+01 lbeta0 = 1.182415579e-05 wbeta0 = 1.031701894e-04 pbeta0 = -1.251454397e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -7.302708231e-01 lkt1 = 5.168481685e-08 wkt1 = 3.971856586e-07 pkt1 = -4.817862039e-14   kt2 = -2.477320583e-01 lkt2 = 2.751982327e-08 wkt2 = 1.898301259e-07 pkt2 = -2.302639427e-14   at = 1.343166196e+05 lat = -7.312039154e-03 wat = -6.026717928e-02 pat = 7.310408846e-9   ute = -3.209663455e+00 lute = 1.759048271e-07 wute = 1.143960347e-06 pute = -1.387623901e-13   ua1 = -2.511895887e-09 lua1 = 2.757580690e-16 wua1 = 1.908460677e-15 pua1 = -2.314962801e-22   ub1 = 2.190926994e-19 lub1 = 2.715631657e-26 wub1 = 4.365759719e-25 pub1 = -5.295666539e-32   uc1 = 6.038902328e-10 luc1 = -7.195567343e-17 wuc1 = -5.272229302e-16 puc1 = 6.395214144e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.64 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.65 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.66 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.170316381e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.387112143e-8   k1 = 6.063790645e-01 lk1 = -2.881841689e-7   k2 = -8.594952435e-02 lk2 = 1.142071145e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.537690438e+05 lvsat = -6.038822173e-1   ua = -8.520891125e-10 lua = -5.004191656e-16   ub = 2.204410149e-18 lub = 7.012749237e-25   uc = -5.909317978e-12 luc = 1.113807635e-16   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214003729e-02 lu0 = 5.030387991e-10   a0 = 2.008729703e+00 la0 = -3.240761624e-7   keta = 1.759108995e-01 lketa = -6.933176282e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.281942499e-01 lags = 3.611563944e-06 pags = 8.077935669e-28   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.036281567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.603596488e-8   nfactor = {1.749350581e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.555897014e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 7.131267544e-01 ldsub = -6.035184771e-7   voffl = 0.0   minv = 0.0   pclm = 1.664834555e-01 lpclm = 1.320987568e-7   pdiblc1 = 0.39   pdiblc2 = 3.512850715e-03 lpdiblc2 = 1.598689531e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.853776267e-05 lalpha0 = 3.163787912e-10   alpha1 = 0.0   beta0 = 1.449521854e+01 lbeta0 = 1.299897675e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470596215e-01 lkt1 = -4.166103278e-8   kt2 = -3.566027875e-02 lkt2 = -2.773576563e-9   at = 6.702214770e+04 lat = -3.465249173e-2   ute = -1.240106715e+00 lute = 2.337455558e-7   ua1 = 1.883327245e-09 lua1 = 3.163790093e-16   ub1 = -1.050270605e-18 lub1 = -1.638514265e-24   uc1 = 1.338950523e-10 luc1 = -2.777712061e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.67 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.260063464e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.448520205e-9   k1 = 4.583535850e-01 lk1 = -8.223055605e-10   k2 = -2.203242067e-02 lk2 = -9.875158843e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.730062600e+03 lvsat = 7.564845687e-2   ua = -7.352140101e-10 lua = -7.273088020e-16   ub = 2.383451972e-18 lub = 3.537010318e-25   uc = 5.799009160e-11 luc = -1.266716032e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.687039536e-02 lu0 = -8.680005323e-9   a0 = 2.227453906e+00 la0 = -7.486854573e-7   keta = -2.459161360e-01 lketa = 1.255751958e-7   a1 = 0.0   a2 = 0.38689047   ags = 1.236107797e+00 lags = 3.806543807e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.188184317e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.452915869e-9   nfactor = {1.005735986e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.879893114e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.470650000e-05 lcit = -9.136728450e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 5.626152760e-04 leta0 = -1.215550353e-10   etab = -5.264411170e-04 letab = 5.133014043e-11   dsub = 2.417621702e-01 ldsub = 3.115415901e-7   voffl = 0.0   minv = 0.0   pclm = 2.558127930e-01 lpclm = -4.131628605e-8   pdiblc1 = 0.39   pdiblc2 = 8.975871500e-03 lpdiblc2 = 5.381533057e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.972691479e-04 lalpha0 = -1.413931643e-10 walpha0 = 1.033975766e-25   alpha1 = 0.0   beta0 = 2.158497514e+01 lbeta0 = -7.643677381e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.675692870e-01 lkt1 = -1.845619147e-9   kt2 = -5.062018750e-02 lkt2 = 2.626809429e-8   at = 2.151566470e+04 lat = 5.368924372e-2   ute = -1.144926840e+00 lute = 4.897286449e-8   ua1 = 2.094023910e-09 lua1 = -9.264642648e-17   ub1 = -2.053097310e-18 lub1 = 3.082732179e-25   uc1 = 2.918378297e-11 luc1 = -7.449521901e-17 puc1 = -5.877471754e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.68 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.438365440e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.033504477e-8   k1 = 4.438791340e-01 lk1 = 1.280249517e-8   k2 = -2.170477869e-02 lk2 = -1.018356824e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.611888860e+04 lvsat = 5.457385496e-2   ua = -1.212585306e-09 lua = -2.779592013e-16   ub = 2.725777112e-18 lub = 3.147037747e-26   uc = 3.374147540e-11 luc = 1.015806211e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214094266e-02 lu0 = -4.228171494e-9   a0 = 1.832745096e+00 la0 = -3.771460549e-7   keta = -2.118113260e-01 lketa = 9.347233816e-8   a1 = 0.0   a2 = 0.38689047   ags = 2.888505226e+00 lags = -1.174747319e-6   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.083733401e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.379048837e-9   nfactor = {1.050183549e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.461508205e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 5.0e-6   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.575917150e-03 leta0 = 1.891445537e-9   etab = -7.780927660e-04 letab = 2.882098376e-10   dsub = 1.956246419e-01 ldsub = 3.549708455e-7   voffl = 0.0   minv = 0.0   pclm = 1.122479820e-01 lpclm = 9.382127054e-8   pdiblc1 = 0.39   pdiblc2 = 2.117781524e-02 lpdiblc2 = -6.104156585e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.571117306e-05 lalpha0 = 7.791121185e-11 palpha0 = 1.232595164e-32   alpha1 = 0.0   beta0 = 1.767369287e+01 lbeta0 = 2.917322269e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.685150100e-01 lkt1 = -9.554100870e-10   kt2 = -1.116694420e-02 lkt2 = -1.086924362e-8   at = 7.604376820e+04 lat = 2.361939893e-3   ute = -1.060861620e+00 lute = -3.015772709e-8   ua1 = 2.467526220e-09 lua1 = -4.442241509e-16   ub1 = -2.108207100e-18 lub1 = 3.601480632e-25   uc1 = -8.371733260e-11 luc1 = 3.177860108e-17 wuc1 = -4.930380658e-32   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.69 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.900716256e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.073858628e-8   k1 = 3.752351760e-01 lk1 = 4.309507383e-8   k2 = -2.572775116e-02 lk2 = -8.408230486e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.591013100e+05 lvsat = -4.111287603e-3   ua = -1.581778528e-09 lua = -1.150342324e-16   ub = 2.641693184e-18 lub = 6.857661490e-26   uc = 6.818598102e-11 luc = -5.042298220e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.448039904e-02 lu0 = -8.475735971e-10   a0 = 5.675289840e-01 la0 = 1.811938154e-7   keta = 2.074182187e-02 lketa = -9.153365992e-9   a1 = 0.0   a2 = 0.38689047   ags = 3.998001480e-01 lags = -7.648176831e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.314017785e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.783401020e-9   nfactor = {2.693661497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.911599775e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.174000000e-06 lcit = 1.688413800e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.588613096e-03 leta0 = 5.363834004e-11   etab = 6.365430149e-03 letab = -2.864226825e-09 wetab = -3.101927297e-25 petab = 2.711709362e-31   dsub = 1.497870141e+00 ldsub = -2.197100933e-7   voffl = 0.0   minv = 0.0   pclm = 1.458467640e-01 lpclm = 7.899412805e-8   pdiblc1 = 0.39   pdiblc2 = 3.543015120e-03 lpdiblc2 = 1.678080708e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.346591437e-04 lalpha0 = 4.304869513e-10 palpha0 = -7.395570986e-32   alpha1 = 0.0   beta0 = 1.996294063e+01 lbeta0 = 1.907077232e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702591400e-01 lkt1 = -1.857255180e-10   kt2 = -4.445217720e-02 lkt2 = 3.819529698e-09 wkt2 = -2.646977960e-23   at = 1.030174912e+05 lat = -9.541564067e-3   ute = -1.212683320e+00 lute = 3.684118912e-8   ua1 = 1.707830040e-09 lua1 = -1.089702267e-16   ub1 = -1.623408644e-18 lub1 = 1.462065046e-25   uc1 = -2.619246032e-11 luc1 = 6.392874939e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.70 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.146155529e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.456383956e-8   k1 = 3.755851429e-01 lk1 = 4.302812517e-8   k2 = -4.657930326e-02 lk2 = -4.419328570e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.439678529e+05 lvsat = -1.216257252e-3   ua = -2.066109318e-09 lua = -2.238175224e-17   ub = 3.773712230e-18 lub = -1.479786286e-25   uc = 6.084055744e-11 luc = -3.637118691e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.314101586e-02 lu0 = -2.504349593e-9   a0 = 4.139458714e+00 la0 = -5.021163420e-7   keta = 1.042213333e-01 lketa = -2.512299653e-08 pketa = -3.155443621e-30   a1 = 0.0   a2 = 0.38689047   ags = -1.896612143e+00 lags = 3.628219029e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.525896395e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.836638845e-9   nfactor = {8.020766929e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.827441752e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.866428571e-05 lcit = -1.657477857e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.210286556e-01 leta0 = 2.370162185e-08 weta0 = 2.646977960e-23 peta0 = -3.944304526e-30   etab = 1.111025482e-02 letab = -3.771911785e-9   dsub = 3.674835515e-01 ldsub = -3.467138701e-9   voffl = 0.0   minv = 0.0   pclm = 1.105167186e+00 lpclm = -1.045238686e-7   pdiblc1 = -6.670428571e-01 lpdiblc1 = 2.022122986e-07 ppdiblc1 = 5.048709793e-29   pdiblc2 = 8.696794286e-03 lpdiblc2 = 6.921627531e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.050656864e-03 lalpha0 = -3.127740010e-10   alpha1 = 0.0   beta0 = 3.268607917e+01 lbeta0 = -5.268591715e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.141323571e-01 lkt1 = -1.092277908e-8   kt2 = -3.077280571e-02 lkt2 = 1.202665933e-9   at = 1.693021714e+04 lat = 6.926931461e-3   ute = 2.611745714e-01 lute = -2.451078255e-7   ua1 = 3.523893743e-09 lua1 = -4.563832130e-16   ub1 = -3.115483286e-18 lub1 = 4.316403836e-25 wub1 = -7.346839693e-40   uc1 = 1.229221143e-12 luc1 = 1.147107275e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.71 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.684310663e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.683166134e-08 wvth0 = 3.418216171e-08 pvth0 = -4.146296216e-15   k1 = 7.674691000e-01 lk1 = -4.507398830e-9   k2 = -1.420406273e-01 lk2 = 7.160130031e-09 wk2 = -8.224025046e-09 pk2 = 9.975742381e-16   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.491298222e+04 lvsat = 9.586098556e-03 wvsat = 8.125032152e-02 pvsat = -9.855664000e-9   ua = -7.686647969e-10 lua = -1.797617726e-16 wua = -1.268217426e-15 pua = 1.538347738e-22   ub = 1.942735858e-18 lub = 7.411880530e-26 wub = 4.424220881e-25 pub = -5.366579929e-32   uc = 1.099604169e-10 luc = -9.595357643e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.644080706e-02 lu0 = -1.691614266e-09 wu0 = -9.994051836e-09 pu0 = 1.212278488e-15   a0 = 0.0   keta = 3.564042735e-01 lketa = -5.571278718e-08 wketa = -3.787281987e-07 pketa = 4.593973050e-14   a1 = 0.0   a2 = 0.38689047   ags = 6.422606667e-01 lags = 5.485663113e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.043695168e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.987537952e-09 wvoff = 1.573733188e-12 pvoff = -1.908938357e-19   nfactor = {3.572517613e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.331030835e-08 wnfactor = -2.309292695e-06 pnfactor = 2.801172040e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.021666667e-05 lcit = 1.845781667e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.119086574e-01 leta0 = -1.668367422e-8   etab = -7.449575150e-02 letab = 6.612096782e-9   dsub = 5.789025160e-01 ldsub = -2.911225910e-8   voffl = 0.0   minv = 0.0   pclm = -1.824672185e-01 lpclm = 5.166618460e-08 wpclm = 1.385900517e-07 ppclm = -1.681097327e-14   pdiblc1 = 1.0   pdiblc2 = -5.810851194e-03 lpdiblc2 = 2.451940150e-09 wpdiblc2 = 5.948034576e-09 ppdiblc2 = -7.214965940e-16   pdiblcb = 0.0   drout = -2.078783057e+01 ldrout = 2.945458829e-06 wdrout = 2.069712970e-05 pdrout = -2.510561833e-12   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.860635655e-03 lalpha0 = -1.684244284e-10 walpha0 = 2.148315020e-11 palpha0 = -2.605906119e-18   alpha1 = 0.0   beta0 = 4.611887097e+01 lbeta0 = -2.156256817e-06 wbeta0 = 4.932722841e-06 pbeta0 = -5.983392807e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.032541950e-01 lkt1 = 1.201769985e-08 wkt1 = 1.184530356e-07 pkt1 = -1.436835322e-14   kt2 = -2.501823667e-02 lkt2 = 5.046367077e-10   at = 1.086564168e+05 lat = -4.199456554e-03 wat = -3.839570541e-02 pat = 4.657399066e-9   ute = -1.867538333e+00 lute = 1.310504983e-8   ua1 = -2.728383667e-10 lua1 = 4.160391877e-18   ub1 = 7.312954000e-19 lub1 = -3.497387102e-26   uc1 = -1.466192333e-11 luc1 = 3.074703100e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.72 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.73 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.4230883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.53326   k2 = -0.056972508   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 200550.0   ua = -9.7905716e-10   ub = 2.38234e-18   uc = 2.2350587e-11   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 0.03226767   a0 = 1.926504   keta = 0.0   a1 = 0.0   a2 = 0.38689047   ags = 0.488144   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5576398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 0.08   etab = -0.07   dsub = 0.56   voffl = 0.0   minv = 0.0   pclm = 0.2   pdiblc1 = 0.39   pdiblc2 = 0.0075691   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.1734937e-5   alpha1 = 0.0   beta0 = 17.793363   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -0.25763   kt2 = -0.036364   at = 58230.0   ute = -1.1808   ua1 = 1.9636e-9   ub1 = -1.466e-18   uc1 = 6.3418e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.74 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.170316381e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.387112143e-8   k1 = 6.063790645e-01 lk1 = -2.881841689e-7   k2 = -8.594952435e-02 lk2 = 1.142071145e-7   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.537690438e+05 lvsat = -6.038822173e-01 wvsat = 2.220446049e-16   ua = -8.520891125e-10 lua = -5.004191656e-16   ub = 2.204410149e-18 lub = 7.012749237e-25   uc = -5.909317978e-12 luc = 1.113807635e-16 puc = 4.701977403e-38   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 3.214003729e-02 lu0 = 5.030387991e-10   a0 = 2.008729703e+00 la0 = -3.240761624e-7   keta = 1.759108995e-01 lketa = -6.933176282e-7   a1 = 0.0   a2 = 0.38689047   ags = -4.281942499e-01 lags = 3.611563944e-06 pags = 1.615587134e-27   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.036281567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.603596488e-8   nfactor = {1.749350581e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.555897014e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 1.571666750e-01 leta0 = -3.041370162e-7   etab = -1.374601750e-01 letab = 2.658807877e-7   dsub = 7.131267544e-01 ldsub = -6.035184771e-7   voffl = 0.0   minv = 0.0   pclm = 1.664834555e-01 lpclm = 1.320987568e-7   pdiblc1 = 0.39   pdiblc2 = 3.512850715e-03 lpdiblc2 = 1.598689531e-8   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -3.853776267e-05 lalpha0 = 3.163787912e-10 palpha0 = 9.860761315e-32   alpha1 = 0.0   beta0 = 1.449521854e+01 lbeta0 = 1.299897675e-5   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.470596215e-01 lkt1 = -4.166103278e-8   kt2 = -3.566027875e-02 lkt2 = -2.773576563e-9   at = 6.702214770e+04 lat = -3.465249173e-2   ute = -1.240106715e+00 lute = 2.337455558e-7   ua1 = 1.883327245e-09 lua1 = 3.163790093e-16   ub1 = -1.050270605e-18 lub1 = -1.638514265e-24   uc1 = 1.338950523e-10 luc1 = -2.777712061e-16   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.75 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {2.343911281e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.784311436e-07 wvth0 = 1.250001877e-07 pvth0 = -2.426628644e-13   k1 = 5.889829475e-01 lk1 = -2.544130869e-07 wk1 = -8.521606460e-08 pk1 = 1.654299462e-13   k2 = -6.109242333e-02 lk2 = 6.595202432e-08 wk2 = 2.548079273e-08 pk2 = -4.946586293e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.822403500e+04 lvsat = -1.072769175e-02 wvsat = -2.902564290e-02 pvsat = 5.634748055e-8   ua = 1.160305674e-09 lua = -4.407081166e-15 wua = -1.236542266e-15 pua = 2.400499501e-21   ub = 2.861387226e-18 lub = -5.741146770e-25 wub = -3.117810630e-25 pub = 6.052605776e-31   uc = -5.577096778e-11 luc = 2.081771842e-16 wuc = 7.421202708e-17 puc = -1.440678082e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 7.330840028e-02 lu0 = -7.941710427e-08 wu0 = -2.377033251e-08 pu0 = 4.614534650e-14   a0 = 2.978646259e+00 la0 = -2.206975173e-06 wa0 = -4.900403319e-07 pa0 = 9.513152963e-13   keta = -3.487845534e-01 lketa = 3.252736544e-07 wketa = 6.710621206e-08 pketa = -1.302732895e-13   a1 = 0.0   a2 = 0.38689047   ags = 1.931307736e+00 lags = -9.689372607e-07 wags = -4.535136801e-07 pags = 8.804061073e-13   b0 = 1.126553268e-06 lb0 = -2.186977859e-12 wb0 = -7.349070245e-13 pb0 = 1.426675007e-18   b1 = 1.122083285e-08 lb1 = -2.178300282e-14 wb1 = -7.319910313e-15 pb1 = 1.421014189e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.070810629e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.747971620e-07 wvoff = 5.757812753e-08 pvoff = -1.117764190e-13   nfactor = {-4.332284519e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.105068852e-05 wnfactor = 3.482257677e-06 pnfactor = -6.760106828e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 4.411428083e-05 lcit = -6.622605338e-11 wcit = -1.918416583e-11 pcit = 3.724222112e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.609631626e-03 leta0 = 4.095427876e-09 weta0 = 1.417065267e-09 peta0 = -2.750948802e-15   etab = 2.249124054e-03 letab = -5.336874525e-09 wetab = -1.810639939e-09 petab = 3.514995314e-15   dsub = -1.597586712e+00 ldsub = 3.882269575e-06 wdsub = 1.199899243e-06 pdsub = -2.329364401e-12   voffl = 0.0   minv = 0.0   pclm = 4.461399506e-01 lpclm = -4.107983970e-07 wpclm = -1.241599212e-07 ppclm = 2.410316551e-13   pdiblc1 = 0.39   pdiblc2 = -9.892160683e-03 lpdiblc2 = 4.201004393e-08 wpdiblc2 = 1.230856079e-08 ppdiblc2 = -2.389460907e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.404700603e-04 lalpha0 = -6.135190955e-10 walpha0 = -1.586521152e-10 palpha0 = 3.079913512e-16   alpha1 = 0.0   beta0 = 2.821975280e+01 lbeta0 = -1.364446160e-05 wbeta0 = -4.328197205e-06 pbeta0 = 8.402329233e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.852863162e-01 lkt1 = -1.615815503e-07 wkt1 = -5.367729598e-08 pkt1 = 1.042037347e-13   kt2 = -1.037776921e-01 lkt2 = 1.294627580e-07 wkt2 = 3.467729815e-08 pkt2 = -6.731903890e-14   at = 5.968108267e+04 lat = -2.040128218e-02 wat = -2.489721041e-02 pat = 4.833295457e-8   ute = -9.302500399e-01 lute = -3.677792075e-07 wute = -1.400444105e-07 pute = 2.718682142e-13   ua1 = 2.755110823e-09 lua1 = -1.376014451e-15 wua1 = -4.312600478e-16 pua1 = 8.372051308e-22   ub1 = -3.058255259e-18 lub1 = 2.259586344e-24 wub1 = 6.557147880e-25 pub1 = -1.272939118e-30   uc1 = 5.455079542e-10 luc1 = -1.076835333e-15 wuc1 = -3.368240731e-16 puc1 = 6.538765731e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.76 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {8.270669807e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.794546365e-07 wvth0 = -2.500003754e-07 pvth0 = 1.103251657e-13   k1 = 1.826204091e-01 lk1 = 1.280959705e-07 wk1 = 1.704321292e-07 pk1 = -7.521169862e-14   k2 = 5.641522662e-02 lk2 = -4.465792658e-08 wk2 = -5.096158547e-08 pk2 = 2.248934767e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -6.286905620e+04 lvsat = 9.384423500e-02 wvsat = 5.805128579e-02 pvsat = -2.561803242e-8   ua = -5.003624675e-09 lua = 1.395026472e-15 wua = 2.473084532e-15 pua = -1.091372204e-21   ub = 1.769906604e-18 lub = 4.532960327e-25 wub = 6.235621260e-25 pub = -2.751779662e-31   uc = 2.612635941e-10 luc = -9.024744889e-17 wuc = -1.484240542e-16 puc = 6.549953510e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -4.073506718e-02 lu0 = 2.793201165e-08 wu0 = 4.754066502e-08 pu0 = -2.097969547e-14   a0 = 3.303603888e-01 la0 = 2.858563164e-07 wa0 = 9.800806638e-07 pa0 = -4.325095969e-13   keta = -6.074491290e-03 lketa = 2.680673006e-09 wketa = -1.342124241e-07 pketa = 5.922794277e-14   a1 = 0.0   a2 = 0.38689047   ags = 1.498105348e+00 lags = -5.611638532e-07 wags = 9.070273603e-07 pags = -4.002711741e-13   b0 = -2.253106536e-06 lb0 = 9.942959145e-13 wb0 = 1.469814049e-12 pb0 = -6.486289398e-19   b1 = -2.244166571e-08 lb1 = 9.903507078e-15 wb1 = 1.463982063e-14 pb1 = -6.460552842e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {6.815192252e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.427964722e-08 wvoff = -1.151562551e-07 pvoff = 5.081845535e-14   nfactor = {1.172622456e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.065186078e-06 wnfactor = -6.964515353e-06 pnfactor = 3.073440625e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -5.381556167e-05 lcit = 2.595530736e-11 wcit = 3.836833165e-11 pcit = -1.693194476e-17   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.768576654e-03 leta0 = -2.577957837e-11 weta0 = -2.834130533e-09 peta0 = 1.250701804e-15   etab = -6.329223107e-03 letab = 2.737923657e-09 wetab = 3.621279878e-09 petab = -1.598070810e-15   dsub = 3.874322406e+00 ldsub = -1.268438478e-06 wdsub = -2.399798487e-06 pdsub = 1.059031072e-12   voffl = 0.0   minv = 0.0   pclm = -2.684063331e-01 lpclm = 2.618040198e-07 wpclm = 2.483198425e-07 ppclm = -1.095835465e-13   pdiblc1 = 0.39   pdiblc2 = 5.891387961e-02 lpdiblc2 = -2.275708179e-08 wpdiblc2 = -2.461712159e-08 ppdiblc2 = 1.086353576e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -5.221129978e-04 lalpha0 = 2.925603371e-10 walpha0 = 3.173042304e-10 palpha0 = -1.400263569e-16   alpha1 = 0.0   beta0 = 4.404137551e+00 lbeta0 = 8.773177029e-06 wbeta0 = 8.656394409e-06 pbeta0 = -3.820066853e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -4.330809515e-01 lkt1 = 7.166753992e-08 wkt1 = 1.073545920e-07 pkt1 = -4.737558143e-14   kt2 = 9.514806507e-02 lkt2 = -5.778605721e-08 wkt2 = -6.935459630e-08 pkt2 = 3.060618335e-14   at = -2.870677310e+02 lat = 3.604673779e-02 wat = 4.979442082e-02 pat = -2.197427791e-8   ute = -1.490215220e+00 lute = 1.593160167e-07 wute = 2.800888211e-07 pute = -1.236031967e-13   ua1 = 1.145352394e-09 lua1 = 1.392511586e-16 wua1 = 8.625200956e-16 pua1 = -3.806301182e-22   ub1 = -9.789120223e-20 lub1 = -5.270043425e-25 wub1 = -1.311429576e-24 pub1 = 5.787338718e-31   uc1 = -1.116365675e-09 luc1 = 4.874863146e-16 wuc1 = 6.736481462e-16 puc1 = -2.972809269e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.77 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.900716256e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.073858628e-8   k1 = 3.752351760e-01 lk1 = 4.309507383e-8   k2 = -2.572775116e-02 lk2 = -8.408230486e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.591013100e+05 lvsat = -4.111287603e-3   ua = -1.581778528e-09 lua = -1.150342324e-16   ub = 2.641693184e-18 lub = 6.857661490e-26   uc = 6.818598102e-11 luc = -5.042298220e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.448039904e-02 lu0 = -8.475735971e-10   a0 = 5.675289840e-01 la0 = 1.811938154e-7   keta = 2.074182187e-02 lketa = -9.153365992e-9   a1 = 0.0   a2 = 0.38689047   ags = 3.998001480e-01 lags = -7.648176831e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.314017785e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.783401020e-9   nfactor = {2.693661497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.911599775e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.174000000e-06 lcit = 1.688413800e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.588613096e-03 leta0 = 5.363834004e-11   etab = 6.365430149e-03 letab = -2.864226825e-09 wetab = -1.033975766e-25 petab = 4.930380658e-32   dsub = 1.497870141e+00 ldsub = -2.197100933e-7   voffl = 0.0   minv = 0.0   pclm = 1.458467640e-01 lpclm = 7.899412805e-8   pdiblc1 = 0.39   pdiblc2 = 3.543015120e-03 lpdiblc2 = 1.678080708e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.346591437e-04 lalpha0 = 4.304869513e-10 palpha0 = 7.395570986e-32   alpha1 = 0.0   beta0 = 1.996294063e+01 lbeta0 = 1.907077232e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702591400e-01 lkt1 = -1.857255180e-10   kt2 = -4.445217720e-02 lkt2 = 3.819529698e-9   at = 1.030174912e+05 lat = -9.541564067e-3   ute = -1.212683320e+00 lute = 3.684118912e-8   ua1 = 1.707830040e-09 lua1 = -1.089702267e-16   ub1 = -1.623408644e-18 lub1 = 1.462065046e-25   uc1 = -2.619246032e-11 luc1 = 6.392874939e-18 wuc1 = 1.232595164e-32   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.78 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {9.496174452e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.186497016e-07 wvth0 = -2.185384845e-07 pvth0 = 4.180641208e-14   k1 = -4.744407283e-02 lk1 = 1.239536141e-07 wk1 = 2.759631089e-07 pk1 = -5.279174272e-14   k2 = 1.431838883e-02 lk2 = -1.606905707e-08 wk2 = -3.972660943e-08 pk2 = 7.599700385e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.281597235e+04 lvsat = 1.430809749e-02 wvsat = 5.293942925e-02 pvsat = -1.012731282e-8   ua = 3.247438635e-09 lua = -1.038863476e-15 wua = -3.466293007e-15 pua = 6.631018522e-22   ub = 7.817739437e-18 lub = -9.216010333e-25 wub = -2.638121148e-24 pub = 5.046725757e-31   uc = -2.021312397e-10 luc = 4.666938611e-17 wuc = 1.715496519e-16 puc = -3.281744841e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 1.035758675e-01 lu0 = -1.597853671e-08 wu0 = -4.594817547e-08 pu0 = 8.789885968e-15   a0 = 4.139458714e+00 la0 = -5.021163420e-7   keta = 1.218294596e+00 lketa = -2.382452117e-07 wketa = -7.267656931e-07 pketa = 1.390302771e-13   a1 = 0.0   a2 = 0.38689047   ags = -1.843557545e+00 lags = 3.526725583e-07 wags = -3.461016722e-08 pags = 6.620924990e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-5.239093750e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.887010425e-08 wvoff = 2.422304294e-07 pvoff = -4.633868115e-14   nfactor = {-1.759738214e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.728193670e-07 wnfactor = 1.671199955e-06 pnfactor = -3.197005514e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 7.280163095e-05 lcit = -1.201395200e-11 wcit = -3.531649717e-11 pcit = 6.756045908e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.392987320e-01 leta0 = 2.719668746e-08 weta0 = 1.191848432e-08 peta0 = -2.280006051e-15   etab = -1.125005278e-01 letab = 1.987483093e-08 wetab = 8.063749403e-08 petab = -1.542595261e-14   dsub = 1.422137270e-01 ldsub = 3.962697873e-08 wdsub = 1.469547700e-07 pdsub = -2.811244751e-14   voffl = 0.0   minv = 0.0   pclm = 1.838403390e+00 lpclm = -2.447919544e-07 wpclm = -4.783266376e-07 ppclm = 9.150388578e-14   pdiblc1 = -1.107224061e+01 lpdiblc1 = 2.192726629e-06 wpdiblc1 = 6.787830755e-06 ppdiblc1 = -1.298512023e-12   pdiblc2 = -1.360779195e-02 lpdiblc2 = 4.959030100e-09 wpdiblc2 = 1.455039683e-08 ppdiblc2 = -2.783490914e-15   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.400864096e-03 lalpha0 = -3.797686445e-10 walpha0 = -2.284576878e-10 palpha0 = 4.370395567e-17   alpha1 = 0.0   beta0 = 3.543371185e+01 lbeta0 = -1.052481304e-06 wbeta0 = -1.792418181e-06 pbeta0 = 3.428895980e-13   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = 1.661283558e-01 lkt1 = -8.366665347e-08 wkt1 = -2.480630761e-07 pkt1 = 4.745446646e-14   kt2 = -1.292702916e-01 lkt2 = 2.004523499e-08 wkt2 = 6.425483494e-08 pkt2 = -1.229194992e-14   at = -2.969286458e+04 lat = 1.584592699e-02 wat = 3.041456736e-02 pat = -5.818306736e-9   ute = 4.539035205e-01 lute = -2.819768735e-07 wute = -1.257267299e-07 pute = 2.405152343e-14   ua1 = 5.216010606e-09 lua1 = -7.800851689e-16 wua1 = -1.103852435e-15 pua1 = 2.111669709e-22   ub1 = -5.877787189e-18 lub1 = 9.600691203e-25 wub1 = 1.801988951e-24 pub1 = -3.447204864e-31   uc1 = -1.768350038e-10 luc1 = 3.521079351e-17 wuc1 = 1.161601972e-16 puc1 = -2.222144572e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.79 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-5.019613663e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.742680827e-08 wvth0 = 6.672176651e-07 pvth0 = -6.563580887e-14   k1 = 1.754537270e+00 lk1 = -9.462672275e-08 wk1 = -6.439139207e-07 pk1 = 5.878934096e-14   k2 = -3.044053618e-01 lk2 = 2.259213388e-08 wk2 = 9.769460951e-08 pk2 = -9.069493473e-15   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.034984284e+05 lvsat = -1.488668443e-02 wvsat = -8.091439432e-02 pvsat = 6.109155984e-9   ua = -1.683188784e-08 lua = 1.396758826e-15 wua = 9.210626126e-15 pua = -8.746084386e-22   ub = -7.381704805e-18 lub = 9.220915533e-25 wub = 6.525220955e-24 pub = -6.068408214e-31   uc = 1.172686932e-09 luc = -1.200960582e-16 wuc = -6.932696424e-16 puc = 7.208513199e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = -1.830991156e-01 lu0 = 1.879513874e-08 wu0 = 1.266993167e-07 pu0 = -1.215225484e-14   a0 = 0.0   keta = -2.822747071e+00 lketa = 2.519331424e-07 wketa = 1.695191181e-06 pketa = -1.547530917e-13   a1 = 0.0   a2 = 0.38689047   ags = 5.184666039e-01 lags = 6.615902906e-08 wags = 8.075705685e-08 pags = -7.373119291e-15   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {7.620646276e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.711854227e-08 wvoff = -5.652167403e-07 pvoff = 5.160466054e-14   nfactor = {7.483847539e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.484275848e-07 wnfactor = -4.860848773e-06 pnfactor = 4.726369593e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -1.365371389e-04 lcit = 1.337884078e-11 wcit = 8.240516005e-11 pcit = -7.523591113e-18   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.545388356e-01 leta0 = -2.057580949e-08 weta0 = -2.780979676e-08 peta0 = 2.539034444e-15   etab = 2.139294079e-01 letab = -1.972112027e-08 wetab = -1.881541527e-07 petab = 1.717847414e-14   dsub = 1.104532107e+00 ldsub = -7.710224071e-08 wdsub = -3.428944634e-07 pdsub = 3.130626451e-14   voffl = 0.0   minv = 0.0   pclm = -6.801048018e-01 lpclm = 6.070308919e-08 wpclm = 4.632239292e-07 ppclm = -2.270619798e-14   pdiblc1 = 2.527879476e+01 lpdiblc1 = -2.216653962e-06 wpdiblc1 = -1.583827176e-05 ppdiblc1 = 1.446034212e-12   pdiblc2 = -6.499971085e-02 lpdiblc2 = 1.119286986e-08 wpdiblc2 = 4.455988717e-08 ppdiblc2 = -6.423642092e-15   pdiblcb = 0.0   drout = 5.745555683e+01 ldrout = -6.545464063e-06 wdrout = -3.034494407e-05 pdrout = 3.680841716e-12   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 1.034995354e-03 lalpha0 = -9.278876604e-11 walpha0 = 5.600896010e-10 palpha0 = -5.194683045e-17   alpha1 = 0.0   beta0 = 2.724559836e+01 lbeta0 = -5.926313646e-08 wbeta0 = 1.724470223e-05 pbeta0 = -1.966313108e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -8.427295747e-01 lkt1 = 3.870781350e-08 wkt1 = 4.051447996e-07 pkt1 = -3.177964886e-14   kt2 = 2.048092305e-01 lkt2 = -2.047861104e-08 wkt2 = -1.499279482e-07 pkt2 = 1.368842167e-14   at = 2.139409646e+05 lat = -1.370685649e-02 wat = -1.070780802e-01 pat = 1.085955141e-8   ute = -2.317239214e+00 lute = 5.416274028e-08 wute = 2.933623698e-07 pute = -2.678398436e-14   ua1 = -6.295540426e-09 lua1 = 6.162659713e-16 wua1 = 3.928909688e-15 pua1 = -3.993070747e-22   ub1 = 7.176671175e-18 lub1 = -6.234366792e-25 wub1 = -4.204640887e-24 pub1 = 3.838837129e-31   uc1 = 4.008212683e-10 luc1 = -3.485891229e-17 wuc1 = -2.710404600e-16 puc1 = 2.474599400e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.80 nmos  lmin = 8e-06 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.989500939e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.266087979e-8   k1 = 7.114214577e-01 wk1 = -1.001890957e-7   k2 = -1.161978331e-01 wk2 = 3.330536155e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.626896858e+05 wvsat = -2.036492523e-1   ua = -2.921559758e-10 wua = -3.862788809e-16   ub = 8.587053423e-19 wub = 8.568159498e-25   uc = 1.290402884e-11 wuc = 5.312271980e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.702382988e-02 wu0 = 2.948873491e-9   a0 = 3.146076880e+00 wa0 = -6.858268091e-7   keta = 4.323500000e-01 wketa = -2.431320225e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.737432051e+00 wags = 2.376252692e-6   b0 = -6.370178385e-07 wb0 = 3.582269815e-13   b1 = -6.344902538e-09 wb1 = 3.568055943e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-4.397552128e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -3.726050612e-8   nfactor = {3.980787014e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.362656836e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.458481970e-01 weta0 = -1.494997336e-7   etab = -3.028038462e-01 wetab = 1.309172429e-7   dsub = 1.557730769e+00 wdsub = -5.610738981e-7   voffl = 0.0   minv = 0.0   pclm = 5.273493846e-02 wpclm = 8.281450736e-8   pdiblc1 = 0.39   pdiblc2 = -5.454279731e-03 wpdiblc2 = 7.323697592e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.134901703e-04 walpha0 = 8.729083908e-11   alpha1 = 0.0   beta0 = 4.132290300e+00 wbeta0 = 7.682304233e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.645808577e-01 wkt1 = 3.908814823e-9   kt2 = -5.170244769e-02 wkt2 = 8.625576060e-9   at = -3.094052462e+04 wat = 5.014504452e-2   ute = -1.594525692e+00 wute = 2.326586431e-7   ua1 = 1.483358923e-09 wua1 = 2.700635696e-16   ub1 = -3.425634615e-20 wub1 = -8.051410437e-25   uc1 = 1.485177831e-10 wuc1 = -4.785586301e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.81 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.989500939e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.266087979e-8   k1 = 7.114214577e-01 wk1 = -1.001890957e-7   k2 = -1.161978331e-01 wk2 = 3.330536155e-8   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.626896858e+05 wvsat = -2.036492523e-1   ua = -2.921559758e-10 wua = -3.862788809e-16   ub = 8.587053423e-19 wub = 8.568159498e-25   uc = 1.290402884e-11 wuc = 5.312271980e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.702382988e-02 wu0 = 2.948873491e-9   a0 = 3.146076880e+00 wa0 = -6.858268091e-7   keta = 4.323500000e-01 wketa = -2.431320225e-7   a1 = 0.0   a2 = 0.38689047   ags = -3.737432051e+00 wags = 2.376252692e-6   b0 = -6.370178385e-07 wb0 = 3.582269815e-13   b1 = -6.344902538e-09 wb1 = 3.568055943e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-4.397552128e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -3.726050612e-8   nfactor = {3.980787014e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.362656836e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.458481970e-01 weta0 = -1.494997336e-7   etab = -3.028038462e-01 wetab = 1.309172429e-7   dsub = 1.557730769e+00 wdsub = -5.610738981e-7   voffl = 0.0   minv = 0.0   pclm = 5.273493846e-02 wpclm = 8.281450736e-8   pdiblc1 = 0.39   pdiblc2 = -5.454279731e-03 wpdiblc2 = 7.323697592e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -1.134901703e-04 walpha0 = 8.729083908e-11   alpha1 = 0.0   beta0 = 4.132290300e+00 wbeta0 = 7.682304233e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.645808577e-01 wkt1 = 3.908814823e-9   kt2 = -5.170244769e-02 wkt2 = 8.625576060e-9   at = -3.094052462e+04 wat = 5.014504452e-2   ute = -1.594525692e+00 wute = 2.326586431e-7   ua1 = 1.483358923e-09 wua1 = 2.700635696e-16   ub1 = -3.425634615e-20 wub1 = -8.051410437e-25   uc1 = 1.485177831e-10 wuc1 = -4.785586301e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.82 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.727503723e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.032609626e-07 wvth0 = -3.133343018e-08 pvth0 = -4.464487717e-14   k1 = 1.027717657e+00 lk1 = -1.246618211e-06 wk1 = -2.369397575e-07 pk1 = 5.389753834e-13   k2 = -2.415457188e-01 lk2 = 4.940336219e-07 wk2 = 8.749951994e-08 pk2 = -2.135954364e-13   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.225479911e+06 lvsat = -2.612255115e+00 wvsat = -4.902066062e-01 pvsat = 1.129408499e-6   ua = 2.570784974e-10 lua = -2.164697829e-15 wua = -6.237404054e-16 pua = 9.359071065e-22   ub = 8.902186545e-20 lub = 3.033553487e-24 wub = 1.189588601e-24 pub = -1.311556850e-30   uc = -1.093417986e-10 luc = 4.818074796e-16 wuc = 5.816525547e-17 puc = -2.083094638e-22   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.647172023e-02 lu0 = 2.176029759e-09 wu0 = 3.187578098e-09 pu0 = -9.408064664e-16   a0 = 3.501766295e+00 la0 = -1.401878692e-06 wa0 = -8.396091277e-07 pa0 = 6.061022525e-13   keta = 1.193299956e+00 lketa = -2.999132063e-06 wketa = -5.721287362e-07 pketa = 1.296674748e-12   a1 = 0.0   a2 = 0.38689047   ags = -7.701299857e+00 lags = 1.562279219e-05 wags = 4.090030938e-06 pags = -6.754514201e-12   b0 = -6.370178385e-07 wb0 = 3.582269815e-13   b1 = -6.344902538e-09 wb1 = 3.568055943e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.539977831e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.126255758e-07 wvoff = -4.961522859e-08 pvoff = 4.869366769e-14   nfactor = {4.810083612e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.268506681e-06 wnfactor = -1.721203220e-06 pnfactor = 1.413138864e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 6.796534254e-01 leta0 = -1.315626547e-06 weta0 = -2.938204241e-07 peta0 = 5.688111374e-13   etab = -5.946209955e-01 letab = 1.150138931e-06 wetab = 2.570843874e-07 petab = -4.972625666e-13   dsub = 2.220121772e+00 ldsub = -2.610681658e-06 wdsub = -8.474586480e-07 pdsub = 1.128728215e-12   voffl = 0.0   minv = 0.0   pclm = -9.224989846e-02 lpclm = 5.714287378e-07 wpclm = 1.454987016e-07 ppclm = -2.470572148e-13   pdiblc1 = 0.39   pdiblc2 = -2.300067808e-02 lpdiblc2 = 6.915561981e-08 wpdiblc2 = 1.490988292e-08 ppdiblc2 = -2.989943223e-14   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -4.607313446e-04 lalpha0 = 1.368581640e-09 walpha0 = 2.374205608e-10 palpha0 = -5.917062722e-16   alpha1 = 0.0   beta0 = -1.013472151e+01 lbeta0 = 5.623057365e-05 wbeta0 = 1.385064679e-05 pbeta0 = -2.431128852e-11   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.188558396e-01 lkt1 = -1.802160137e-07 wkt1 = -1.586039674e-08 pkt1 = 7.791639354e-14   kt2 = -4.865831196e-02 lkt2 = -1.199785215e-08 wkt2 = 7.309443977e-09 pkt2 = 5.187271379e-15   at = 7.092277378e+03 lat = -1.498986825e-01 wat = 3.370156258e-02 pat = 6.480869538e-8   ute = -1.851072855e+00 lute = 1.011129333e-06 wute = 3.435768090e-07 pute = -4.371617672e-13   ua1 = 1.136117509e-09 lua1 = 1.368582584e-15 wua1 = 4.201933948e-16 pua1 = -5.917066800e-22   ub1 = 1.764093079e-18 lub1 = -7.087834590e-24 wub1 = -1.582657418e-24 pub1 = 3.064425285e-30   uc1 = 4.533852472e-10 luc1 = -1.201574137e-15 wuc1 = -1.796653111e-16 puc1 = 5.195005779e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.83 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {6.442295790e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.296316213e-07 wvth0 = -1.054724652e-07 pvth0 = 9.928123146e-14   k1 = 2.969578800e-01 lk1 = 1.720057445e-07 wk1 = 7.900423207e-08 pk1 = -7.436668365e-14   k2 = 6.198646193e-02 lk2 = -9.521340046e-08 wk2 = -4.373261839e-08 pk2 = 4.116551369e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3.195114628e+05 lvsat = 3.870366392e-01 wvsat = 1.777704143e-01 pvsat = -1.673352910e-7   ua = -5.496296392e-10 lua = -5.986353237e-16 wua = -2.749601426e-16 pua = 2.588199822e-22   ub = 5.326372237e-19 lub = 2.172362992e-24 wub = 9.977915008e-25 pub = -9.392211397e-31   uc = 2.458299577e-10 luc = -2.076874509e-16 wuc = -9.539325338e-17 puc = 8.979366940e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.170784653e-02 lu0 = 1.142413779e-08 wu0 = 5.247238895e-09 pu0 = -4.939225972e-15   a0 = 3.927860477e+00 la0 = -2.229055327e-06 wa0 = -1.023830947e-06 pa0 = 9.637320706e-13   keta = -5.602098578e-01 lketa = 4.049565392e-07 wketa = 1.860012320e-07 pketa = -1.750829597e-13   a1 = 0.0   a2 = 0.38689047   ags = -9.832055374e-01 lags = 2.580955682e-06 wags = 1.185462859e-06 pags = -1.115876189e-12   b0 = -1.416939332e-06 lb0 = 1.514061595e-12 wb0 = 6.954260391e-13 pb0 = -6.546045306e-19   b1 = -1.411317144e-08 lb1 = 1.508054041e-14 wb1 = 6.926667001e-15 pb1 = -6.520071648e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.000450369e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.036864224e-07 wvoff = -4.762437557e-08 pvoff = 4.482882473e-14   nfactor = {5.288931136e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.198093380e-06 wnfactor = -1.928232947e-06 pnfactor = 1.815045673e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 3.724265645e-03 leta0 = -3.445268739e-09 weta0 = -1.582451864e-09 peta0 = 1.489561939e-15   etab = -4.198807904e-03 letab = 3.952337880e-09 wetab = 1.815354597e-09 petab = -1.708793282e-15   dsub = 1.454502737e+00 ldsub = -1.124385426e-06 wdsub = -5.164432584e-07 pdsub = 4.861280391e-13   voffl = 0.0   minv = 0.0   pclm = 1.624032459e-01 lpclm = 7.707058866e-08 wpclm = 3.539941465e-08 ppclm = -3.332146901e-14   pdiblc1 = 0.39   pdiblc2 = 1.369357296e-02 lpdiblc2 = -2.078929725e-09 wpdiblc2 = -9.548765181e-10 ppdiblc2 = 8.988252665e-16   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.909450711e-04 lalpha0 = -2.847777855e-10 walpha0 = -1.308017375e-10 palpha0 = 1.231236755e-16   alpha1 = 0.0   beta0 = 1.594062183e+01 lbeta0 = 5.610509619e-06 wbeta0 = 2.576972096e-06 pbeta0 = -2.425703834e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -3.645410532e-01 lkt1 = 1.026026914e-07 wkt1 = 4.712660534e-08 pkt1 = -4.436027361e-14   kt2 = -7.657007557e-02 lkt2 = 4.218725453e-08 wkt2 = 1.937709497e-08 pkt2 = -1.823965950e-14   at = -2.161804790e+05 lat = 2.835407195e-01 wat = 1.302335388e-01 pat = -1.225888301e-7   ute = -1.587969081e+00 lute = 5.003659756e-07 wute = 2.298238920e-07 pute = -2.163332295e-13   ua1 = 1.589867105e-09 lua1 = 4.877184944e-16 wua1 = 2.240147573e-16 pua1 = -2.108650910e-22   ub1 = -1.878025245e-18 lub1 = -1.739028667e-26 wub1 = -7.987560228e-27 pub1 = 7.518690442e-33   uc1 = -3.570267350e-10 luc1 = 3.716786447e-16 wuc1 = 1.707163094e-16 puc1 = -1.606952620e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.84 nmos  lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {3.825033186e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.673130760e-8   k1 = 4.856916800e-01 lk1 = -5.649381384e-9   k2 = -3.420731355e-02 lk2 = -4.666199603e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.036075760e+04 lvsat = 4.828891817e-2   ua = -6.058572126e-10 lua = -5.457083088e-16   ub = 2.878757188e-18 lub = -3.603973006e-26   uc = -2.671773805e-12 luc = 2.622722898e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.380421444e-02 lu0 = -9.375173330e-09 wu0 = -1.323488980e-23   a0 = 2.073190768e+00 la0 = -4.832547299e-7   keta = -2.447380000e-01 lketa = 1.080028794e-7   a1 = 0.0   a2 = 0.38689047   ags = 3.111028546e+00 lags = -1.272946860e-6   b0 = 3.605932040e-07 lb0 = -1.591297809e-13   b1 = 3.591624280e-09 lb1 = -1.584983795e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.366249158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.088371549e-9   nfactor = {-6.584386451e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.400165795e-06 pnfactor = 2.019483917e-28   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.441300000e-05 lcit = -4.153956900e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -2.271221573e-03 leta0 = 2.198283379e-09 weta0 = 1.550963649e-25 peta0 = -3.328006944e-31   etab = 1.103250000e-04 letab = -1.038489225e-10   dsub = -3.931240000e-01 ldsub = 6.147856212e-07 pdsub = -5.048709793e-29   voffl = 0.0   minv = 0.0   pclm = 1.731689180e-01 lpclm = 6.693686149e-8   pdiblc1 = 0.39   pdiblc2 = 1.513843444e-02 lpdiblc2 = -3.438977838e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 4.213387759e-05 lalpha0 = 4.355819100e-11   alpha1 = 0.0   beta0 = 1.979738803e+01 lbeta0 = 1.980135591e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.421774360e-01 lkt1 = -1.257818149e-8   kt2 = -2.818188300e-02 lkt2 = -3.360551132e-9   at = 8.825995960e+04 lat = -3.029065371e-3   ute = -9.921467200e-01 lute = -6.048161246e-8   ua1 = 2.679130460e-09 lua1 = -5.376051020e-16   ub1 = -2.429943440e-18 lub1 = 5.021303101e-25   uc1 = 8.155047360e-11 luc1 = -4.115408180e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.85 nmos  lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {4.900716256e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.073858628e-8   k1 = 3.752351760e-01 lk1 = 4.309507383e-8   k2 = -2.572775116e-02 lk2 = -8.408230486e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.591013100e+05 lvsat = -4.111287603e-3   ua = -1.581778528e-09 lua = -1.150342324e-16   ub = 2.641693184e-18 lub = 6.857661490e-26   uc = 6.818598102e-11 luc = -5.042298220e-18   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.448039904e-02 lu0 = -8.475735971e-10   a0 = 5.675289840e-01 la0 = 1.811938154e-7   keta = 2.074182187e-02 lketa = -9.153365992e-9   a1 = 0.0   a2 = 0.38689047   ags = 3.998001480e-01 lags = -7.648176831e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.314017785e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.783401020e-9   nfactor = {2.693661497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.911599775e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.174000000e-06 lcit = 1.688413800e-12   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.588613096e-03 leta0 = 5.363834004e-11   etab = 6.365430149e-03 letab = -2.864226825e-09 wetab = -7.237830360e-25 petab = -3.204747427e-31   dsub = 1.497870141e+00 ldsub = -2.197100933e-7   voffl = 0.0   minv = 0.0   pclm = 1.458467640e-01 lpclm = 7.899412805e-8   pdiblc1 = 0.39   pdiblc2 = 3.543015120e-03 lpdiblc2 = 1.678080708e-9   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = -8.346591437e-04 lalpha0 = 4.304869513e-10 walpha0 = 5.169878828e-26 palpha0 = -2.465190329e-32   alpha1 = 0.0   beta0 = 1.996294063e+01 lbeta0 = 1.907077232e-6   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.702591400e-01 lkt1 = -1.857255180e-10   kt2 = -4.445217720e-02 lkt2 = 3.819529698e-9   at = 1.030174912e+05 lat = -9.541564067e-3   ute = -1.212683320e+00 lute = 3.684118912e-8   ua1 = 1.707830040e-09 lua1 = -1.089702267e-16   ub1 = -1.623408644e-18 lub1 = 1.462065046e-25   uc1 = -2.619246032e-11 luc1 = 6.392874939e-18 wuc1 = -6.162975822e-33 puc1 = -1.469367939e-39   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.25e-6   sbref = 1.24e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.86 nmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {5.610009529e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.430736658e-8   k1 = 4.432878714e-01 lk1 = 3.007659320e-8   k2 = -5.632553299e-02 lk2 = -2.554874822e-9   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.569556171e+05 lvsat = -3.700816559e-3   ua = -2.916503762e-09 lua = 1.402987049e-16   ub = 3.126495286e-18 lub = -2.416602716e-26   uc = 1.029272681e-10 luc = -1.168830644e-17   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 2.186843357e-02 lu0 = -3.479046022e-10   a0 = 4.139458714e+00 la0 = -5.021163420e-7   keta = -7.407793525e-02 lketa = 8.985653546e-9   a1 = 0.0   a2 = 0.38689047   ags = -1.905103143e+00 lags = 3.644462312e-7   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-9.316263466e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.531747188e-9   nfactor = {1.212076411e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.043112291e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = -1.181046637e-01 leta0 = 2.314226219e-08 weta0 = -3.308722450e-24 peta0 = 1.577721810e-30   etab = 3.089325550e-02 letab = -7.556399815e-9   dsub = 4.035363375e-01 ldsub = -1.036403666e-8   voffl = 0.0   minv = 0.0   pclm = 9.878181000e-01 lpclm = -8.207498853e-8   pdiblc1 = 9.982328571e-01 lpdiblc1 = -1.163549456e-7   pdiblc2 = 1.226648000e-02 lpdiblc2 = 9.281876000e-12   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 2.994608761e-03 lalpha0 = -3.020519989e-10   alpha1 = 0.0   beta0 = 3.224634068e+01 lbeta0 = -4.427371978e-7   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -2.749903000e-01 lkt1 = 7.193453900e-10   kt2 = -1.500900429e-02 lkt2 = -1.812949280e-9   at = 2.439190000e+04 lat = 5.499511530e-3   ute = 2.303297143e-01 lute = -2.392072043e-7   ua1 = 3.253082829e-09 lua1 = -4.045770851e-16   ub1 = -2.673396771e-18 lub1 = 3.470692334e-25   uc1 = 2.972709657e-11 luc1 = -4.304536294e-18   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.1e-6   sbref = 1.1e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_01v8_lvt__model.87 nmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.148e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.935e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = -6.175e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -1.33e-8   dwb = -1.08e-8   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = -3.0e-7   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 0.0   xn = 0.0   rnoia = 0.912   rnoib = 0.26   tnoia = 25000000.0   tnoib = 9900000.0   epsrox = 3.9   toxe = {3.932304e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(3.932304e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {9.033449613e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -8.583369481e-08 wvth0 = -1.230563482e-07 pvth0 = 1.492673504e-14   k1 = 6.094960667e-01 lk1 = 9.915539113e-9   k2 = 3.614158715e-02 lk2 = -1.377113650e-08 wk2 = -9.381196721e-08 pk2 = 1.137939162e-14   k3 = 1.65   dvt0 = 0.07665   dvt1 = 0.1252   dvt2 = -0.05637   dvt0w = 0.0   dvt1w = 5300000.0   dvt2w = -0.032   w0 = 1.0e-7   k3b = 1.6   vfb = 0.0   phin = 0.0   lpe0 = 2.3802e-7   lpeb = -4.9152e-8   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.289240880e+05 lvsat = -3.005920756e-04 wvsat = 1.725748602e-02 pvsat = -2.093333054e-9   ua = -1.456835607e-09 lua = -3.675904233e-17 wua = 5.644655025e-16 pua = -6.846966545e-23   ub = 7.708208101e-18 lub = -5.799277917e-25 wub = -1.960591568e-24 pub = 2.378197572e-31   uc = -2.991750540e-10 luc = 3.708670523e-17 wuc = 1.344319457e-16 puc = -1.630659501e-23   rdsw = 103.65   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = 4.021634726e-02 lu0 = -2.573506532e-09 wu0 = 1.117866179e-09 pu0 = -1.355971675e-16   a0 = 0.0   keta = -5.000693549e-01 lketa = 6.065841275e-08 wketa = 3.890333672e-07 pketa = -4.718974745e-14   a1 = 0.0   a2 = 0.38689047   ags = 6.620730000e-01 lags = 5.304776510e-8   b0 = 0.0   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.430413979e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.464854679e-08 wvoff = 4.633111352e-12 pvoff = -5.619964070e-19   nfactor = {-7.712940909e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.286915830e-06 wnfactor = 3.685065211e-06 pnfactor = -4.469984101e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = 1.0e-5   cdsc = 3.8556e-37   cdscb = -0.00011484   cdscd = 4.7984e-6   eta0 = 2.050860095e-01 leta0 = -1.606076646e-8   etab = -1.206560864e-01 letab = 1.082653536e-8   dsub = 4.947793487e-01 ldsub = -2.143181392e-8   voffl = 0.0   minv = 0.0   pclm = 1.436240667e-01 lpclm = 2.032574771e-8   pdiblc1 = -2.885643333e+00 lpdiblc1 = 3.547592363e-07 wpdiblc1 = 5.293955920e-23 ppdiblc1 = -1.262177448e-29   pdiblc2 = 1.423899667e-02 lpdiblc2 = -2.299843957e-10   pdiblcb = 0.0   drout = 3.4946   pscbe1 = 450000000.0   pscbe2 = 1.0e-8   pvag = 0.0   delta = 0.01   alpha0 = 3.286611766e-03 lalpha0 = -3.374719633e-10 walpha0 = -7.061068882e-10 palpha0 = 8.565076554e-17   alpha1 = 0.0   beta0 = 1.325499095e+02 lbeta0 = -1.260956009e-05 wbeta0 = -4.197317711e-05 pbeta0 = 5.091346384e-12   fprout = 0.0   pdits = 1.4427e-15   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.148e-9   kt1 = -1.222800333e-01 lkt1 = -1.780440996e-8   kt2 = -6.180044000e-02 lkt2 = 3.862851872e-9   at = -8.201705655e+04 lat = 1.840691796e-02 wat = 5.935391300e-02 pat = -7.199629647e-9   ute = -1.795567000e+00 lute = 6.534067100e-9   ua1 = 1.795197183e-09 lua1 = -2.277355563e-16 wua1 = -6.209166062e-16 pua1 = 7.531718433e-23   ub1 = -3.002398000e-19 lub1 = 5.920529274e-26   uc1 = -8.115696600e-11 luc1 = 9.145700496e-18 wuc1 = -6.162975822e-33 puc1 = -7.346839693e-40   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 9.0e+41   noib = 1.0e+27   noic = 800000000000.0   em = 41000000.0   af = 1.0   ef = 1.2   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.2928   jss = 0.00275   jsws = 6.0e-10   xtis = 2.0   bvs = 11.9   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0012287   tpbsw = 0.0   tpbswg = 0.0   tcj = 0.000792   tcjsw = 1.0e-5   tcjswg = 0.0   cgdo = 2.228188563e-10   cgso = 2.228188563e-10   cgbo = 1.0e-14   capmod = 2.0   xpart = 0.0   cgsl = 2.151675e-11   cgdl = 2.151675e-11   cf = 1.0e-14   clc = 1.0e-7   cle = 0.6   dlc = 2.4805e-8   dwc = -6.175e-9   vfbcv = -1.0   acde = 0.38008   moin = 23.81   noff = 3.8661   voffcv = -0.16994   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099678423   mjs = 0.42197   pbs = 0.7477   cjsws = 2.7168e-11   mjsws = 0.001   pbsws = 0.1   cjswgs = 1.5099e-10   mjswgs = 0.8   pbswgs = 0.79644   saref = 1.04e-6   sbref = 1.04e-6   wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54













* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__nfet_01v8_lvt





















