** Translated using xdm 2.6.0 on Nov_14_2022_16_05_13_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__RF_PFET_01V8_B__TOXE_MULT=1.0365 SKY130_FD_PR__RF_PFET_01V8_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_PFET_01V8_B__OVERLAP_MULT=1.1043 SKY130_FD_PR__RF_PFET_01V8_B__AJUNCTION_MULT=1.0625 
+ SKY130_FD_PR__RF_PFET_01V8_B__PJUNCTION_MULT=1.0675 SKY130_FD_PR__RF_PFET_01V8_B__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__RF_PFET_01V8_B__WINT_DIFF=2.252e-8 SKY130_FD_PR__RF_PFET_01V8_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__DLC_DIFF=-1.21275e-8 SKY130_FD_PR__RF_PFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_B__XGW_DIFF=4.504e-8 SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT=1.1125 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT=1.315 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT=1.315 
+ SKY130_FD_PR__RF_PFET_01V8__AW_CAP_MULT_2=1.1125 SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_DIST_MULT_2=1.21 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RGATE_STUB_MULT_2=1.21 SKY130_FD_PR__RF_PFET_01V8__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_PFET_01V8__AW_RS_MULT=1.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_0=-0.025683 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_0=-0.00046629 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_0=0.036263 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_0=-4705.4 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_1=-0.0096007 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_1=-0.00041939 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_1=0.036542 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_1=-19320.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_2=-0.00361 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_2=-0.000495 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_2=0.022214 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_2=-19622.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_3=-0.02462 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_3=-0.0008663 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_3=0.054438 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_3=-17486.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_4=-0.018152 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_4=-0.00068712 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_4=0.046452 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_4=-11488.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_5=-0.016536 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_5=-0.00054677 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_5=0.022396 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_5=-14168.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_6=-0.025252 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_6=-0.0012477 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_6=0.074957 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_6=-15388.0 SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_7=-0.0006238 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_7=-19606.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_7=-0.013565 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_7=0.045593 SKY130_FD_PR__RF_PFET_01V8_BM02__VTH0_DIFF_8=0.026563 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__U0_DIFF_8=-0.0006639 SKY130_FD_PR__RF_PFET_01V8_BM02__VSAT_DIFF_8=-20194.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__B1_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UB_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM02__K2_DIFF_8=-0.013354 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_0=-0.024438 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_0=-0.00066296 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_0=0.049452 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_0=-8761.9 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_1=-0.0094416 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_1=-0.00051496 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_1=0.050655 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_1=-10144.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_2=-0.00053393 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_2=0.029231 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_2=-14879.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_2=-0.0049051 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_3=-0.022453 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_3=-0.00092315 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_3=0.053737 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_3=-16685.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_4=-0.00093397 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_4=0.059286 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_4=-15584.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_4=-0.014614 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_5=0.029916 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_5=-0.00065774 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_5=-21301.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_5=-0.0167 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_5=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_6=0.078414 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_6=-0.0011357 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_6=-13899.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_6=-0.024399 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_7=-0.010627 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_7=0.049986 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_7=-0.00088539 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_7=-18591.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_7=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__K2_DIFF_8=-0.012274 SKY130_FD_PR__RF_PFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_PFET_01V8_BM04__VTH0_DIFF_8=0.038873 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__U0_DIFF_8=-0.000789 SKY130_FD_PR__RF_PFET_01V8_BM04__UA_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__VSAT_DIFF_8=-17257.0 SKY130_FD_PR__RF_PFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_PFET_01V8_BM04__UB_DIFF_8=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_pfet_01v8_b.pm3.spice














