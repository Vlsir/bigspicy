** Translated using xdm 2.6.0 on Nov_14_2022_16_05_03_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_05V0_NVT__TOXE_SLOPE=0.105e-2
.PARAM SKY130_FD_PR__NFET_05V0_NVT__TOXE_SLOPE1=1.205e-2
.PARAM SKY130_FD_PR__NFET_05V0_NVT__TOXE_SLOPE2=2.525e-2
* .param sky130_fd_pr__nfet_05v0_nvt__vth0_slope=0.0012  ; All devices; HSpice Parser Retained (as a comment). Continuing.
.PARAM SKY130_FD_PR__NFET_05V0_NVT__VOFF_SLOPE=0.0035
.PARAM SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_SLOPE=0.02
* .param sky130_fd_pr__nfet_05v0_nvt__lint_slope=0.0e-9  ; All devices; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__nfet_05v0_nvt__wint_slope=0.0e-9  ; All devices; HSpice Parser Retained (as a comment). Continuing.
