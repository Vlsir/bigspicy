** Translated using xdm 2.6.0 on Nov_14_2022_16_05_16_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_B__TOXE_MULT=1.052 SKY130_FD_PR__RF_NFET_01V8_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_NFET_01V8_B__OVERLAP_MULT=0.9600 SKY130_FD_PR__RF_NFET_01V8_B__AJUNCTION_MULT=1.2169 
+ SKY130_FD_PR__RF_NFET_01V8_B__PJUNCTION_MULT=1.2474 SKY130_FD_PR__RF_NFET_01V8_B__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__RF_NFET_01V8_B__WINT_DIFF=3.2175e-8 SKY130_FD_PR__RF_NFET_01V8_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__DLC_DIFF=-17.422e-9 SKY130_FD_PR__RF_NFET_01V8_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_B__XGW_DIFF=6.4250e-8 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_0=0.032714 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_0=20474.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_0=0.0083532 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_0=0.00017601 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_1=0.032194 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_1=21175.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_1=0.014272 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_1=-0.00050746 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_2=0.018697 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_2=32392.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_2=0.031744 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_2=-0.0018379 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_3=0.036104 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_3=12645.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_3=0.0022323 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_3=-0.0069942 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_4=0.0098858 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_4=23380.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_4=0.0131 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_4=-0.0040868 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_5=0.0085637 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_5=21055.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_5=0.032731 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_5=-0.0019994 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_6=-0.0048122 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_6=0.015103 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_6=4095.2 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_6=0.0010067 SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_7=0.011492 SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_7=-0.0042353 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_7=0.0051454 SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_7=18771.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__K2_DIFF_8=0.030405 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__U0_DIFF_8=-0.0042395 SKY130_FD_PR__RF_NFET_01V8_BM02__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__RDSW_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__KT1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM02__VTH0_DIFF_8=0.0015836 
+ SKY130_FD_PR__RF_NFET_01V8_BM02__VSAT_DIFF_8=20830.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_0=0.0072696 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_0=-0.0014397 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_0=0.057292 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_0=10629.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_1=0.018201 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_1=-0.0021915 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_1=0.020199 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_1=24240.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_2=0.033909 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_2=-0.0024784 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_2=0.01762 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_2=39930.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_3=11859.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_3=0.0020408 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_3=-0.0072915 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_3=0.030316 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_4=27029.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_4=0.015422 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_4=-0.0070125 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_4=0.0054988 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_5=55116.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_5=0.034152 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_5=-0.0062872 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_5=0.0021981 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_6=4091.9 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_6=0.0010631 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_6=-0.0047075 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_6=0.015982 SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_7=-0.0056998 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_7=12177.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_7=0.014379 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_7=-0.0040004 SKY130_FD_PR__RF_NFET_01V8_BM04__VTH0_DIFF_8=-0.0017169 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__U0_DIFF_8=-0.0057354 SKY130_FD_PR__RF_NFET_01V8_BM04__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VOFF_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UB_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__VSAT_DIFF_8=47784.0 SKY130_FD_PR__RF_NFET_01V8_BM04__AGS_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__B0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_BM04__K2_DIFF_8=0.03191
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*





* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*














* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_b.pm3.spice














