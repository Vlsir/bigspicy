** Translated using xdm 2.6.0 on Nov_14_2022_16_05_34_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 05
.PARAM 
+ SKY130_FD_PR__NFET_G5V0D16V0__TOXE_MULT=1.0 SKY130_FD_PR__NFET_G5V0D16V0__TOXP_MULT=1.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__OVERLAP_MULT=1.0 SKY130_FD_PR__NFET_G5V0D16V0__AJUNCTION_MULT=9.9505e-1 
+ SKY130_FD_PR__NFET_G5V0D16V0__PJUNCTION_MULT=1.0144e+0 SKY130_FD_PR__NFET_G5V0D16V0__CJS_MULT=1.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CJSWS_MULT=1.0 SKY130_FD_PR__NFET_G5V0D16V0__CJSWGS_MULT=1.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGDO_MULT=1.0 SKY130_FD_PR__NFET_G5V0D16V0__CGSO_MULT=1.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGDL_MULT=1.0 SKY130_FD_PR__NFET_G5V0D16V0__CGSL_MULT=1.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CF_MULT=1.0 SKY130_FD_PR__NFET_G5V0D16V0__RDIFF_MULT=1.0588 
+ SKY130_FD_PR__NFET_G5V0D16V0__LINT_DIFF=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DLC_DIFF=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__WINT_DIFF=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DWC_DIFF=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_0=1.0521e-2 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_0=-1.4914e-3 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_1=9.8261e-4 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_1=-5.0931e-3 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_2=8.6130e-3 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_2=-1.9057e-3 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_3=1.0853e-2 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_3=-1.3899e-3 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_4=1.7461e-2 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_4=-2.9881e-3 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_4=0.0
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 000, W = 20.0, L = 0.7
* --------------------------------
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 001, W = 5.0, L = 0.7
* --------------------------------
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 002, W = 50.0, L = 0.7
* --------------------------------
*




















* sky130_fd_pr__nfet_g5v0d16v0, Bin 003, W = 20.0, L = 2.2
* --------------------------------
*






















* sky130_fd_pr__nfet_g5v0d16v0, Bin 004, W = 5.0, L = 2.2
* -------------------------------
.INCLUDE sky130_fd_pr__nfet_g5v0d16v0__subcircuit.pm3.spice






















.INCLUDE sky130_fd_pr__nfet_g5v0d16v0.pm3.spice
