** Translated using xdm 2.6.0 on Nov_14_2022_16_05_13_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 2
.PARAM 
+ SKY130_FD_PR__PFET_G5V0D16V0__TOXE_MULT=1.0365 SKY130_FD_PR__PFET_G5V0D16V0__RSHP_MULT=1.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__SOVERLAP_MULT=1.70 SKY130_FD_PR__PFET_G5V0D16V0__DOVERLAP_MULT=1.70 
+ SKY130_FD_PR__PFET_G5V0D16V0__AJUNCTION_MULT=1.0559e+0 SKY130_FD_PR__PFET_G5V0D16V0__PJUNCTION_MULT=1.0542e+0 
+ SKY130_FD_PR__PFET_G5V0D16V0__WINT_DIFF=2.252e-8 SKY130_FD_PR__PFET_G5V0D16V0__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__PFET_G5V0D16V0__DLC_DIFF=-1.21275e-8 SKY130_FD_PR__PFET_G5V0D16V0__DWC_DIFF=2.252e-8 
+ SKY130_FD_PR__PFET_G5V0D16V0__CF_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D16V0__CJSWGS_DIFF=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGC_DIFF=0.0 SKY130_FD_PR__PFET_G5V0D16V0__RDIFF_MULT=1.9011 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGBINV_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__UA_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGBACC_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__NIGBACC_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__DSUB_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__BIGSD_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VSAT_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGSD_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__RDW_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__A0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__LPE0_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGC_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__KETA_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__UB_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__K2_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PDITSD_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VTH0_DIFF_0=-0.105 SKY130_FD_PR__PFET_G5V0D16V0__U0_DIFF_0=-8.94e-3 
+ SKY130_FD_PR__PFET_G5V0D16V0__NIGBINV_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__RDSW_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__B1_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AGIDL_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__B0_DIFF_0=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VOFF_DIFF_0=0.0 SKY130_FD_PR__PFET_G5V0D16V0__JTSSWS_DIFF_0=-4.02e-12 
+ SKY130_FD_PR__PFET_G5V0D16V0__AGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__B0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VOFF_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGBINV_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__CGIDL_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__UA_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__KT1_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AIGBACC_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__NIGBACC_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__DSUB_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__BIGSD_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PCLM_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__AIGSD_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__RDW_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PDITS_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__A0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__ETA0_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__LPE0_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__KETA_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__UB_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__K2_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__PDITSD_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__VTH0_DIFF_1=-0.129 SKY130_FD_PR__PFET_G5V0D16V0__U0_DIFF_1=-6.79e-3 
+ SKY130_FD_PR__PFET_G5V0D16V0__NIGBINV_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__RDSW_DIFF_1=0.0 SKY130_FD_PR__PFET_G5V0D16V0__B1_DIFF_1=0.0 
+ SKY130_FD_PR__PFET_G5V0D16V0__JTSSWS_DIFF_1=-4.02e-12
*
* sky130_fd_pr__pfet_g5v0d16v0__base, Bin 000, W = 27.545, L = 0.66
* ----------------------------------------
*







* sky130_fd_pr__pfet_g5v0d16v0__base, Bin 001, W = 27.545, L = 2.16
* ----------------------------------------
