** Translated using xdm 2.6.0 on Nov_14_2022_16_05_34_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_G5V0D10V5__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_G5V0D10V5__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_G5V0D10V5__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_G5V0D10V5__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__nfet_g5v0d10v5 d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__nfet_g5v0d10v5 d g s b sky130_fd_pr__nfet_g5v0d10v5__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__nfet_g5v0d10v5__model.0 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.1 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.2 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.783366897345+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.2790420190348e-8   k1 = 0.88325   k2 = -0.04100161561805 lk2 = 1.04727100702197e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110468.7325 lvsat = -0.037734056605245   ua = -1.0160370546575e-10 lua = 3.32403078041264e-16   ub = 1.752361942755e-18 lub = -2.79760295671284e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0415573116048 lu0 = 4.32281352469685e-9   a0 = 1.03361118331195 la0 = -7.14172112976905e-7   keta = -0.0172681619955 lketa = -3.17947160955794e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1520662575117 lags = -2.07824090159046e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.012092027505+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.6654862586335e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.259908962315 lpclm = 5.81783684739667e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4994591 lbeta0 = 1.96217094347274e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414270958 lkt1 = 9.05617358525876e-8   kt2 = -0.019151   at = 236939.72 lat = -0.60374490568392   ute = -1.33706986 lute = 3.0187245284196e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.3 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.799231213062+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.82393802725314e-8   k1 = 0.88325   k2 = -0.0425688326357 lk2 = 1.6501771996081e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93779.97715 lvsat = 0.0264673515836301   ua = 1.059936792802e-10 lua = -4.6622115471302e-16 pua = -5.64237288394698e-37   ub = 1.54968606504e-18 lub = 4.99930968436031e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0427638373221 lu0 = -3.18674018396179e-10   a0 = 0.4765335596815 la0 = 1.42889770604271e-6   keta = -0.039268111389 lketa = 5.28387812219236e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.119434808895 lags = 1.04750316972259e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96133159753+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.71273962395545e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60098245601 lpclm = -7.30321270476086e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.859072776 lbeta0 = 1.05443086577469e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577642e-8   kt2 = -0.019151   at = 139103.552 lat = -0.227370537094272   ute = -1.22166028 lute = -1.42106585683921e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.4 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.77849763948+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.00552398633929e-8   k1 = 0.88325   k2 = -0.040704192142 lk2 = 1.3057807109184e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 119885.646358 lvsat = -0.021749453964177   ua = -1.424027673504e-10 lua = -7.43639533655408e-18   ub = 1.763188445e-18 lub = 1.05595061683231e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0411635356998 lu0 = 2.6370606737692e-9   a0 = 1.7025972264586 la0 = -8.35624721603264e-7   keta = 0.003322044888 lketa = -2.58246411595076e-08 pketa = -5.04870979341448e-29   a1 = 0.0   a2 = 0.65972622   ags = 0.152949206474 lags = 4.28496938454126e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.9020982963+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.18708842899521e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.0967492387200001 lpclm = 2.00990422593502e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 27.084637048 lbeta0 = 4.58673660526266e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.38119986 lkt1 = 1.564371284196e-8   kt2 = -0.019151   at = 9224.11200000001 lat = 0.012514970273568   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.0067651972e-18 lub1 = 4.69624259515638e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.5 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78843401736+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.16392669083229e-8   k1 = 0.88325   k2 = -0.036128620909 lk2 = 9.18236233283029e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 85126.2279969999 lvsat = 0.007691286755733   ua = -1.60784842719e-10 lua = 8.13296515159496e-18   ub = 1.6018274894e-18 lub = 2.42265532023053e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.045631465191 lu0 = -1.1472130542643e-9   a0 = -0.59798198177 la0 = 1.11293365965745e-6   keta = -0.08057022444 lketa = 4.52309364695378e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.3435801197 lags = -1.18612020824224e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.8523738453+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.97549704352654e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.9101826875 lpclm = 1.90083366705488e-06 ppclm = 3.23117426778526e-27   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.10834751e-06 lalpha0 = 7.92664763789513e-12   alpha1 = 0.0   beta0 = 22.85343874 lbeta0 = 8.17050233536235e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.33685056 lkt1 = -2.19195233678399e-8   kt2 = -0.019151   at = 7825.35000000001 lat = 0.0136997021049   ute = -1.465198895 lute = 1.4110693168047e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -9.939305129e-18 lub1 = 5.4944025261912e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.6 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7757384111+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.98531464200556e-8   k1 = 0.88325   k2 = -0.012073800896 lk2 = -6.38076944810054e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 83539.70703 lvsat = 0.0087177436100884   ua = -2.9722602282e-10 lua = 9.64084985004205e-17   ub = 1.1918419193e-18 lub = 5.07520456079771e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.037431758785 lu0 = 4.15788219452798e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.8407922064+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.22618122099105e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.031822874 lpclm = -2.60274315776379e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.67118703e-05 lalpha0 = 4.19330842084195e-13   alpha1 = 0.0   beta0 = 32.17877346 lbeta0 = 2.13714132620844e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909599e-8   ua1 = 2.0117e-9   ub1 = -1.670493e-18 lub1 = 1.44596842098e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.7 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.86273265206+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.90320613696912e-8   k1 = 0.88325   k2 = 0.000971042710000009 lk2 = -1.22116319121721e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 102046.556208 lvsat = 0.000445441123410911   ua = 1.47858737334e-10 lua = -1.02538158101775e-16   ub = -9.44912075800003e-19 lub = 1.46261957733354e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.038101135306 lu0 = 3.8586802609123e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.1695064304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.59192468338775e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.128000231999999 lpclm = 4.01393324299248e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.869456438e-05 lalpha0 = -4.93676565395868e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768392001e-8   kt2 = -0.019151   at = -462.432000000059 lat = 0.017370963029952   ute = -1.30083493 lute = 7.75489420979589e-10   ua1 = -1.432830022e-09 lua1 = 1.53965669641369e-15   ub1 = 5.78529723000001e-18 lub1 = -3.18803700964878e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.8 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.9 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.10 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.783366897344999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.27904201903497e-8   k1 = 0.88325   k2 = -0.04100161561805 lk2 = 1.04727100702197e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110468.7325 lvsat = -0.0377340566052449   ua = -1.0160370546575e-10 lua = 3.32403078041264e-16 wua = 7.88860905221012e-31 pua = -3.00926553810506e-36   ub = 1.752361942755e-18 lub = -2.7976029567129e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0415573116048 lu0 = 4.32281352469664e-9   a0 = 1.03361118331195 la0 = -7.14172112976903e-07 wa0 = 1.35525271560688e-20   keta = -0.0172681619955 lketa = -3.17947160955796e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1520662575117 lags = -2.07824090159046e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.012092027505+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.66548625863353e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.259908962315 lpclm = 5.81783684739668e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4994591 lbeta0 = 1.96217094347274e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414270958 lkt1 = 9.05617358525889e-8   kt2 = -0.019151   at = 236939.72 lat = -0.60374490568392   ute = -1.33706986 lute = 3.01872452841955e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.11 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.799231213061999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.82393802725322e-8   k1 = 0.88325   k2 = -0.0425688326357 lk2 = 1.6501771996081e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93779.97715 lvsat = 0.02646735158363   ua = 1.059936792802e-10 lua = -4.66221154713019e-16 wua = -1.97215226305253e-31 pua = -3.76158192263132e-37   ub = 1.54968606504e-18 lub = 4.99930968436029e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0427638373220999 lu0 = -3.18674018396285e-10   a0 = 0.4765335596815 la0 = 1.42889770604271e-6   keta = -0.039268111389 lketa = 5.28387812219235e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.119434808895 lags = 1.04750316972259e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96133159753+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.71273962395545e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60098245601 lpclm = -7.30321270476086e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.859072776 lbeta0 = 1.05443086577468e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577635e-8   kt2 = -0.019151   at = 139103.552 lat = -0.227370537094272   ute = -1.22166028 lute = -1.42106585683916e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.12 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.779602344057306+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.80148659749727e-08 wvth0 = -2.20469294982996e-08 pvth0 = 4.07203701263428e-14   k1 = 0.88325   k2 = -0.0400796286596472 lk2 = 1.19042471011671e-08 wk2 = -1.24646057828678e-08 pk2 = 2.30219523764757e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 127486.824642213 lvsat = -0.0357887238386221 wvsat = -0.151699056180947 pvsat = 2.80186032979422e-7   ua = -1.49239013726612e-10 lua = 5.19005601285932e-18 wua = 1.36433074493939e-16 pua = -2.51989978527262e-22   ub = 1.6593816868986e-18 lub = 2.97324690601902e-25 wub = 2.0717034439111e-24 pub = -3.82640725705565e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0405271650538457 lu0 = 3.81242834765779e-09 wu0 = 1.27002449834683e-08 pu0 = -2.34571746810378e-14   a0 = 1.75957160491531 la0 = -9.40855600971506e-07 wa0 = -1.13705521896909e-06 pa0 = 2.10012507066282e-12   keta = 0.003322044888 lketa = -2.58246411595076e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.0384105981257299 lags = 2.54400899924151e-07 wags = 2.2858822846978e-06 pags = -4.22199257748485e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.903339822086421+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.41639650361122e-08 wnfactor = -2.47775125095605e-08 pnfactor = 4.57637187199855e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.09674923872 lpclm = 2.00990422593502e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 27.1479802003684 lbeta0 = 4.46974268964232e-06 wbeta0 = -1.26415880150749e-06 pbeta0 = 2.33488360816158e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.38119986 lkt1 = 1.56437128419601e-8   kt2 = -0.019151   at = 9224.11200000001 lat = 0.012514970273568   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.0067651972e-18 lub1 = 4.69624259515637e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.13 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.782910494473471+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.5212908886587e-08 wvth0 = 1.10234647491484e-07 pvth0 = -7.13202736419374e-14   k1 = 0.88325   k2 = -0.0392514383207641 lk2 = 1.12027814787979e-08 wk2 = 6.23230289143385e-08 pk2 = -4.03221271851721e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 47120.3365759356 lvsat = 0.0322805664226813 wvsat = 0.758495280904732 pvsat = -4.90735827811429e-7   ua = -1.26603610837942e-10 lua = -1.39818133382031e-17 wua = -6.82165372469693e-16 pua = 4.41351445672674e-22   ub = 2.120861279907e-18 lub = -9.35420639619084e-26 wub = -1.03585172195557e-23 pub = 6.70181562181144e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0488133184207715 lu0 = -3.20582754798129e-09 wu0 = -6.3501224917344e-08 pu0 = 4.10844035043731e-14   a0 = -0.88285387405354 la0 = 1.2972417857584e-06 wa0 = 5.6852760948454e-06 pa0 = -3.67829403949965e-12   keta = -0.08057022444 lketa = 4.52309364695379e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.91627316144135 lags = -4.89136401128293e-07 wags = -1.1429411423489e-05 pags = 7.39466917923744e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.846166216367891+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.57387214229954e-08 wnfactor = 1.23887562547803e-07 pnfactor = -8.01535185425356e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.9101826875 lpclm = 1.90083366705488e-06 ppclm = -6.46234853557053e-27   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.10834751e-06 lalpha0 = 7.92664763789514e-12   alpha1 = 0.0   beta0 = 22.5367229781579 lbeta0 = 8.37541299925358e-06 wbeta0 = 6.32079400753917e-06 pbeta0 = -4.08946523176166e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.33685056 lkt1 = -2.19195233678405e-8   kt2 = -0.019151   at = 7825.34999999998 lat = 0.0136997021049   ute = -1.465198895 lute = 1.41106931680471e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -9.93930512899999e-18 lub1 = 5.49440252619119e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.14 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.775738411099999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.98531464200552e-8   k1 = 0.88325   k2 = -0.012073800896 lk2 = -6.38076944810054e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 83539.7070299999 lvsat = 0.00871774361008848   ua = -2.9722602282e-10 lua = 9.64084985004205e-17   ub = 1.1918419193e-18 lub = 5.07520456079771e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.037431758785 lu0 = 4.157882194528e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.8407922064+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.22618122099107e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.031822874 lpclm = -2.60274315776336e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.67118703e-05 lalpha0 = 4.19330842084195e-13   alpha1 = 0.0   beta0 = 32.1787734599999 lbeta0 = 2.13714132620842e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -1.670493e-18 lub1 = 1.44596842098e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.15 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.895377604079501+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.36238978930782e-08 wvth0 = -6.51505362098337e-07 pvth0 = 2.91213775782881e-13   k1 = 0.88325   k2 = 0.00535553483497164 lk2 = -1.41714385091447e-08 wk2 = -8.75026597616334e-08 pk2 = 3.91124638762137e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123736.609686367 lvsat = -0.00924970912067014 wvsat = -0.43287507780423 pvsat = 1.93489099527402e-7   ua = 9.04067357655688e-11 lua = -7.68579177287086e-17 wua = 1.14658729051767e-15 pua = -5.12508466639332e-22   ub = -2.99298059184676e-18 lub = 2.37807753104722e-24 wub = 4.08739341798481e-23 pub = -1.82700763433136e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0436741320434463 lu0 = 1.3676287412282e-09 wu0 = -1.11222012372209e-07 pu0 = 4.97146824222045e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.47405424987601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.95321079975078e-07 wnfactor = -6.07795463401117e-06 pnfactor = 2.71676063003812e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.00611809398051 lpclm = 1.35531433835597e-06 wpclm = 4.25912567400374e-05 ppclm = -1.90376954852024e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.869456438e-05 lalpha0 = -4.93676565395869e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.440127200000001 lkt1 = 3.10195768391997e-8   kt2 = -0.019151   at = -82837.738590376 lat = 0.0541915718215578 wat = 1.64398936521856 pat = -7.34840230401585e-7   ute = -1.30083493 lute = 7.75489420978319e-10   ua1 = -1.432830022e-09 lua1 = 1.53965669641369e-15   ub1 = 2.1523136984184e-18 lub1 = -1.56414423280125e-24 wub1 = 7.25045712987018e-23 pub1 = -3.24085283065215e-29   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.16 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.17 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.18 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.783366897344999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.27904201903497e-8   k1 = 0.88325   k2 = -0.04100161561805 lk2 = 1.04727100702197e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110468.7325 lvsat = -0.0377340566052453   ua = -1.0160370546575e-10 lua = 3.32403078041264e-16   ub = 1.752361942755e-18 lub = -2.7976029567129e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0415573116048 lu0 = 4.32281352469664e-9   a0 = 1.03361118331195 la0 = -7.14172112976906e-7   keta = -0.0172681619955 lketa = -3.17947160955795e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1520662575117 lags = -2.07824090159046e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.012092027505+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.66548625863353e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.259908962315 lpclm = 5.81783684739669e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4994591 lbeta0 = 1.96217094347273e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414270958 lkt1 = 9.05617358525872e-8   kt2 = -0.019151   at = 236939.72 lat = -0.60374490568392   ute = -1.33706986 lute = 3.01872452841962e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.19 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.799231213062001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.82393802725305e-8   k1 = 0.88325   k2 = -0.0425688326357 lk2 = 1.6501771996081e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93779.97715 lvsat = 0.0264673515836302   ua = 1.059936792802e-10 lua = -4.66221154713019e-16 wua = -9.86076131526265e-32 pua = 3.76158192263132e-37   ub = 1.54968606504e-18 lub = 4.99930968436029e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0427638373221 lu0 = -3.18674018396179e-10   a0 = 0.4765335596815 la0 = 1.4288977060427e-6   keta = -0.039268111389 lketa = 5.28387812219235e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.119434808895 lags = 1.0475031697226e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96133159753+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.71273962395544e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60098245601 lpclm = -7.30321270476086e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.859072776 lbeta0 = 1.05443086577468e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577635e-8   kt2 = -0.019151   at = 139103.552 lat = -0.227370537094272   ute = -1.22166028 lute = -1.42106585683919e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.20 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.770338987826502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.51241552462811e-08 wvth0 = 1.16507942759553e-07 pvth0 = -2.15188539165701e-13   k1 = 0.88325   k2 = -0.0391759692414392 lk2 = 1.02352008069689e-08 wk2 = -2.5980918028105e-08 pk2 = 4.79863918650578e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 124467.791778077 lvsat = -0.0302126124050231 wvsat = -0.106542451769943 pvsat = 1.96782416824761e-7   ua = -1.31344104495032e-10 lua = -2.78615908091391e-17 wua = -1.31226594514844e-16 pua = 2.42373682896592e-22   ub = 1.74833303743661e-18 lub = 1.33032791477108e-25 wub = 7.41230696898164e-25 pub = -1.36904271994115e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0409342713291349 lu0 = 3.06050875668634e-09 wu0 = 6.61103103523484e-09 pu0 = -1.22104817676439e-14   a0 = 2.54892884320106 la0 = -2.39878736908395e-06 wa0 = -1.29437145540385e-05 pa0 = 2.39068595693053e-11   keta = 0.0311667503719283 lketa = -7.72534223624464e-08 wketa = -4.16481836092405e-07 pketa = 7.69236120516966e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.203781496858135 lags = -5.10368348420196e-08 wags = -1.87621181879597e-07 pags = 3.46533696235071e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.89692666609284+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.23189557001504e-08 wnfactor = 7.11460369384894e-08 pnfactor = -1.31405734180871e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.746886340835661 lpclm = -9.99803703094693e-07 wpclm = -9.72430087857138e-06 ppclm = 1.79606475825091e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.25154417103886e-05 lalpha0 = 3.60450083909622e-12 walpha0 = 2.9190058417671e-11 palpha0 = -5.39136292366204e-17   alpha1 = 0.0   beta0 = 27.5273159240528 lbeta0 = 3.76911491869737e-06 wbeta0 = -6.93800005605819e-06 pbeta0 = 1.2814388971539e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.398067260947376 lkt1 = 4.67975662481504e-08 wkt1 = 2.52290911129394e-07 pkt1 = -4.65977780783238e-13   kt2 = -0.019151   at = 9224.11199999999 lat = 0.012514970273568   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.51312457364023e-18 lub1 = 1.40486293876947e-24 wub1 = 7.57377315210441e-24 pub1 = -1.39886529791127e-29   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.21 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.82922727562749+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.47534000851283e-08 wvth0 = -5.82539713797772e-07 pvth0 = 3.76895039271176e-13   k1 = 0.88325   k2 = -0.0437697354118039 lk2 = 1.41260564405414e-08 wk2 = 1.29904590140525e-07 pk2 = -8.4046451156658e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 62215.5008966157 lvsat = 0.0225142064395023 wvsat = 0.532712258849717 pvsat = -3.44657373504143e-7   ua = -2.16078156995841e-10 lua = 4.39069653823111e-17 wua = 6.56132972574215e-16 pua = -4.24508847393901e-22   ub = 1.67610452721695e-18 lub = 1.9420932843401e-25 wub = -3.70615348449081e-24 pub = 2.39782941831678e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0467777870443251 lu0 = -1.88886724485975e-09 wu0 = -3.30551551761733e-08 pu0 = 2.13862226268112e-14   a0 = -4.8296400654823 la0 = 3.85075719660613e-06 wa0 = 6.47185727701923e-05 pa0 = -4.18720105222957e-11   keta = -0.219793751859642 lketa = 1.35306609580662e-07 wketa = 2.08240918046202e-06 pketa = -1.3472895860304e-12   a1 = 0.0   a2 = 0.65972622   ags = 0.0894186677793243 lags = 4.5826880308126e-08 wags = 9.38105909397985e-07 pags = -6.06941389897766e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.878231996335801+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.64848321413152e-08 wnfactor = -3.55730184692447e-07 pnfactor = 2.30152449273436e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -5.1608681980783 lpclm = 4.00398168280189e-06 wpclm = 4.86215043928569e-05 ppclm = -3.14574326411169e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4866138958057e-05 lalpha0 = 1.61349318008252e-12 walpha0 = -1.45950292088355e-10 palpha0 = 9.44277956770762e-17   alpha1 = 0.0   beta0 = 20.6400443597358 lbeta0 = 9.60253751187192e-06 wbeta0 = 3.46900002802918e-05 pbeta0 = -2.24439445213448e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.252513555263119 lkt1 = -7.64843847145351e-08 wkt1 = -1.26145455564697e-06 pkt1 = 8.16143437139815e-13   kt2 = -0.019151   at = 7825.34999999992 lat = 0.0136997021049   ute = -1.465198895 lute = 1.41106931680469e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -7.40750824679887e-18 lub1 = 3.85636538856341e-24 wub1 = -3.78688657605221e-23 pub1 = 2.45006259829371e-29   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.22 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.775738411100001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.98531464200552e-8   k1 = 0.88325   k2 = -0.012073800896 lk2 = -6.38076944810054e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 83539.70703 lvsat = 0.00871774361008837   ua = -2.9722602282e-10 lua = 9.64084985004205e-17   ub = 1.1918419193e-18 lub = 5.07520456079769e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.037431758785 lu0 = 4.157882194528e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.840792206400001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.22618122099103e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.031822874 lpclm = -2.60274315776506e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.67118703e-05 lalpha0 = 4.19330842084208e-13   alpha1 = 0.0   beta0 = 32.17877346 lbeta0 = 2.13714132620842e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909603e-8   ua1 = 2.0117e-9   ub1 = -1.670493e-18 lub1 = 1.44596842098e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.23 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.861044916444746+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.82776671779717e-08 wvth0 = -1.37980778677581e-07 pvth0 = 6.16754763379804e-14   k1 = 0.88325   k2 = 0.00333149231096208 lk2 = -1.32667198375077e-08 wk2 = -5.72284323249251e-08 pk2 = 2.5580308051189e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 87996.9925015471 lvsat = 0.0067253994063034 wvsat = 0.101693384231204 pvsat = -4.54555190439686e-8   ua = 1.62670628352059e-10 lua = -1.09158866020373e-16 wua = 6.57139918226254e-17 pua = -2.93732343488285e-23   ub = -6.41434726177268e-19 lub = 1.32696945073507e-24 wub = 5.70113839090281e-24 pub = -2.54832904479609e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0346170596665455 lu0 = 5.41601329468948e-09 wu0 = 2.42474087473852e-08 pu0 = -1.0838252246359e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.13148089590428+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.4219558677667e-07 wnfactor = -9.53979466062946e-07 pnfactor = 4.26415465617612e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.26211855798051 lpclm = -5.52527689757474e-07 wpclm = -2.12500734802323e-05 ppclm = 9.49848534463512e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.869456438e-05 lalpha0 = -4.93676565395868e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768391999e-8   kt2 = -0.019151   at = 81912.8745903759 lat = -0.0194496457616538 wat = -0.820236299314803 pat = 3.66634142485526e-7   ute = -1.30083493 lute = 7.7548942098086e-10   ua1 = -1.43283002200001e-09 lua1 = 1.53965669641369e-15   ub1 = 6.99974823000001e-18 lub1 = -3.73087960433478e-24 pub1 = -1.12103877145985e-44   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.24 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.25 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78882+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.039667   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.92431e-11   ub = 1.71671e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0421082   a0 = 0.9425989   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1494178   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96538+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.26 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.783366897344999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.27904201903463e-8   k1 = 0.88325   k2 = -0.04100161561805 lk2 = 1.04727100702197e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110468.7325 lvsat = -0.0377340566052453   ua = -1.0160370546575e-10 lua = 3.32403078041264e-16 pua = -1.50463276905253e-36   ub = 1.752361942755e-18 lub = -2.79760295671284e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0415573116048 lu0 = 4.32281352469685e-9   a0 = 1.03361118331195 la0 = -7.14172112976903e-7   keta = -0.0172681619955 lketa = -3.17947160955795e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1520662575117 lags = -2.07824090159046e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.012092027505+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.6654862586335e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.259908962315 lpclm = 5.81783684739666e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4994591 lbeta0 = 1.96217094347275e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414270958 lkt1 = 9.05617358525889e-8   kt2 = -0.019151   at = 236939.72 lat = -0.60374490568392   ute = -1.33706986 lute = 3.01872452841955e-07 wute = 6.7762635780344e-21   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.27 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.799231213062001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.82393802725305e-8   k1 = 0.88325   k2 = -0.0425688326357 lk2 = 1.6501771996081e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93779.9771499999 lvsat = 0.0264673515836302   ua = 1.059936792802e-10 lua = -4.66221154713019e-16 wua = -9.86076131526265e-32   ub = 1.54968606504e-18 lub = 4.99930968436029e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0427638373221 lu0 = -3.18674018396179e-10   a0 = 0.4765335596815 la0 = 1.4288977060427e-6   keta = -0.039268111389 lketa = 5.28387812219235e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.119434808895 lags = 1.04750316972259e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96133159753+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.71273962395544e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60098245601 lpclm = -7.30321270476086e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.859072776 lbeta0 = 1.05443086577468e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577644e-8   kt2 = -0.019151   at = 139103.552 lat = -0.227370537094272   ute = -1.22166028 lute = -1.42106585683921e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.28 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.782039734932+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.35130391528847e-8   k1 = 0.88325   k2 = -0.0417852003738 lk2 = 1.50544141792034e-08 wk2 = -2.11758236813575e-22   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 113767.86648 lvsat = -0.0104500001784292   ua = -1.445230274042e-10 lua = -3.52030470082623e-18   ub = 1.8227739101e-18 lub = -4.45845815995806e-27   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.041598208915 lu0 = 1.83422533071982e-9   a0 = 1.249007764729 la0 = 2.14866395884254e-9   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.1849389360094 lags = -1.62348887502576e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.90407177368+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.55158693821291e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.22971304512 lpclm = 8.03961690374008e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.5446962802e-05 lalpha0 = -1.80997757581477e-12   alpha1 = 0.0   beta0 = 26.830541248 lbeta0 = 5.05604799052144e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 9224.11200000001 lat = 0.012514970273568   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.29 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.770723540100001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.30976977488612e-8   k1 = 0.88325   k2 = -0.0307235797500001 lk2 = 5.68537637353348e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 115715.127387 lvsat = -0.0120993029050055   ua = -1.5018354245e-10 lua = 1.27407229575541e-18   ub = 1.3039001639e-18 lub = 4.35020340638995e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0434580991150001 lu0 = 2.58924369782601e-10   a0 = 1.669965326878 la0 = -3.5439649777549e-7   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.183631472023 lags = -1.51274850582728e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.842506458400003+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.33709092543818e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.2778712683 lpclm = 8.44751031192344e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.08533500000005e-07 lalpha0 = 1.1096758704969e-11   alpha1 = 0.0   beta0 = 24.12391774 lbeta0 = 7.34852020906833e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.379199860000001 lkt1 = 5.47988084196013e-9   kt2 = -0.019151   at = 7825.35000000003 lat = 0.0136997021049   ute = -1.465198895 lute = 1.41106931680469e-7   ua1 = 6.21571501100001e-09 lua1 = -2.71993885590685e-15   ub1 = -1.1210631115e-17 lub1 = 6.31693264056939e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.30 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7757384111+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.98531464200552e-8   k1 = 0.88325   k2 = -0.012073800896 lk2 = -6.38076944810055e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 83539.70703 lvsat = 0.00871774361008848   ua = -2.9722602282e-10 lua = 9.64084985004204e-17   ub = 1.1918419193e-18 lub = 5.07520456079771e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.037431758785 lu0 = 4.15788219452797e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.8407922064+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.22618122099107e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.031822874 lpclm = -2.60274315776506e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.67118703e-05 lalpha0 = 4.19330842084195e-13   alpha1 = 0.0   beta0 = 32.17877346 lbeta0 = 2.13714132620845e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -1.670493e-18 lub1 = 1.44596842098e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.31 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.75208868731985+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.0424241853649e-08 wvth0 = 9.46929953237586e-07 pvth0 = -4.23264432077852e-13   k1 = 0.88325   k2 = -0.00110262350631363 lk2 = -1.12847321448069e-08 wk2 = -1.30765754246381e-08 pk2 = 5.84504614275744e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 101675.677888443 lvsat = 0.000611218539956715 wvsat = -0.03450949920121 pvsat = 1.54252630099524e-8   ua = 1.98141252128225e-10 lua = -1.25013738259587e-16 wua = -2.87477934068784e-16 pua = 1.28498611837669e-22   ub = -5.32864326242839e-19 lub = 1.27844000194998e-24 wub = 4.62006947907257e-24 pub = -2.06510637617271e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.033122060592836 lu0 = 6.08425695065059e-09 wu0 = 3.91335749840272e-08 pu0 = -1.74921601478105e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.21029299646343+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.77423492357203e-07 wnfactor = -1.73873582545741e-06 pnfactor = 7.77190571677904e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.128000232 lpclm = 4.01393324299248e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.869456438e-05 lalpha0 = -4.9367656539587e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768392001e-8   kt2 = -0.019151   at = -77713.2631580164 lat = 0.0519010030459491 wat = 0.769210319096364 pat = -3.43826243691608e-7   ute = -1.30083493 lute = 7.75489420979166e-10   ua1 = -1.432830022e-09 lua1 = 1.53965669641369e-15   ub1 = 8.60914054579202e-18 lub1 = -4.45025543800139e-24 wub1 = -1.60252149811743e-23 pub1 = 7.16304674357515e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.32 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.773930725422+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.03589269135717e-7   k1 = 0.88325   k2 = -0.039005199382 wk2 = -4.60435073401634e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 119218.23738 wvsat = -0.0943288333897736   ua = -3.776291806848e-10 wua = 2.215110026237e-15   ub = 2.15421721754e-18 wub = -3.04387246464878e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0412944578918 wu0 = 5.66145447931683e-9   a0 = 1.2299227366222 wa0 = -1.99900042712233e-6   keta = -0.017029449926 wketa = -2.98506783542409e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1698880119244 wags = -1.42417569183323e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.90891626188+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.92835616932181e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.6534245679 wpclm = -2.22198723624721e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.3789217694e-05 walpha0 = -6.48575397402078e-11   alpha1 = 0.0   beta0 = 26.68933959 wbeta0 = -1.87105638442238e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 179829.232 wat = -0.137958074427456   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.33 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.773930725422+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.03589269135713e-7   k1 = 0.88325   k2 = -0.039005199382 wk2 = -4.60435073401613e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 119218.23738 wvsat = -0.0943288333897732   ua = -3.776291806848e-10 wua = 2.215110026237e-15   ub = 2.15421721754e-18 wub = -3.04387246464878e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0412944578918 wu0 = 5.66145447931683e-9   a0 = 1.2299227366222 wa0 = -1.99900042712233e-6   keta = -0.017029449926 wketa = -2.98506783542408e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1698880119244 wags = -1.42417569183323e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.90891626188+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.92835616932178e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.6534245679 wpclm = -2.22198723624721e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.3789217694e-05 walpha0 = -6.48575397402078e-11   alpha1 = 0.0   beta0 = 26.68933959 wbeta0 = -1.87105638442237e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 179829.232 wat = -0.137958074427456   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.34 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.762108010812788+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.27726760204819e-08 wvth0 = 1.47904621341652e-07 pvth0 = -3.47741948345032e-13   k1 = 0.88325   k2 = -0.0397195406622933 lk2 = 5.60542602568351e-09 wk2 = -8.91979034628553e-09 pk2 = 3.38631942213221e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 142215.64473428 lvsat = -0.180460333545331 wvsat = -0.220873046462854 pvsat = 9.92990668365479e-7   ua = -5.2574203144813e-10 lua = 1.16223946635994e-15 wua = 2.95086096846382e-15 pua = -5.77342734314064e-21   ub = 2.32055109417595e-18 lub = -1.305219601288e-24 wub = -3.95306692869417e-24 pub = 7.13443623064162e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0401955254141624 lu0 = 8.62330776696754e-09 wu0 = 9.47436595841243e-09 pu0 = -2.9919862995704e-14   a0 = 1.5409259695701 la0 = -2.44043801489692e-06 wa0 = -3.52954522095213e-06 pa0 = 1.20101635695554e-11   keta = -0.00293450744429405 lketa = -1.10602816324752e-07 wketa = -9.97236494783415e-08 pketa = 5.48292226189223e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.202417148688517 lags = -2.55255680780112e-07 wags = -3.50306657991598e-07 pags = 1.63130276943129e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.928619418336639+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.54610392871056e-07 wnfactor = 5.80744651547907e-07 pnfactor = -1.47451956390316e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.395513550592924 lpclm = 2.02382414205438e-06 wpclm = -9.43442886862708e-07 ppclm = -1.00327196099993e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.55129271216997e-05 lalpha0 = -9.19957837472276e-11 walpha0 = -1.46422997131218e-10 palpha0 = 6.40043002230856e-16   alpha1 = 0.0   beta0 = 26.8014838328953 lbeta0 = -8.79994303979608e-07 wbeta0 = -3.688781909037e-05 pbeta0 = 1.42636667434937e-10   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414270958 lkt1 = 9.05617358525872e-8   kt2 = -0.019151   at = 275839.646473688 lat = -0.753392378229227 wat = -0.270638769654801 pat = 1.04114355791924e-6   ute = -1.33706986 lute = 3.01872452841962e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.35 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.794535772576738+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.19764694967695e-08 wvth0 = 3.26676256516338e-08 pvth0 = 9.55731607565246e-14   k1 = 0.88325   k2 = -0.0432634050859056 lk2 = 1.9238622849218e-08 wk2 = 4.83235446439469e-09 pk2 = -1.9041114335337e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 73043.8726742042 lvsat = 0.085642505164971 wvsat = 0.14426746555829 pvsat = -4.11699769412692e-7   ua = 1.21573265364366e-10 lua = -1.32797341806358e-15 wua = -1.0839197890006e-16 pua = 5.99547591582695e-21   ub = 1.55831895914198e-18 lub = 1.62707675093776e-24 wub = -6.00617031988865e-26 pub = -7.84190036976555e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0438512315785742 lu0 = -5.44014266763837e-09 wu0 = -7.56533675972225e-09 pu0 = 3.56316348051216e-14   a0 = 0.277442505170145 la0 = 2.42016518388121e-06 wa0 = 1.38513778628029e-06 pa0 = -6.89655315370565e-12   keta = -0.0511014773099234 lketa = 7.46948424107462e-08 wketa = 8.23283713885678e-08 pketa = -1.52059349357485e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.114212514707311 lags = 8.40663112807102e-08 wags = 3.63331091303589e-08 pags = 1.43904998269862e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.943205817120531+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.10724064783106e-07 wnfactor = 1.26106637049043e-07 pnfactor = 2.74466512941796e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.58199022372901 lpclm = -2.54053500882672e-06 wpclm = -6.82517319041362e-06 ppclm = 1.25942145235368e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 8.95080162348575e-06 lalpha0 = 1.01883411746446e-11 walpha0 = 3.83778910945096e-11 palpha0 = -7.0883427561084e-17   alpha1 = 0.0   beta0 = 23.8066283661974 lbeta0 = 1.06411727484306e-05 wbeta0 = 3.64871911875259e-07 pbeta0 = -6.73913313026689e-13   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577644e-8   kt2 = -0.019151   at = 148259.630473688 lat = -0.262593842797451 wat = -0.0637016580136174 pat = 2.45059386555174e-7   ute = -1.22166028 lute = -1.42106585683919e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.36 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.76915514368721+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.49011967333842e-08 wvth0 = 8.9642069744115e-08 pvth0 = -9.6578398400634e-15   k1 = 0.88325   k2 = -0.0405000056852206 lk2 = 1.41346628437445e-08 wk2 = -8.94149528841101e-09 pk2 = 6.39899332419866e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 125778.021544817 lvsat = -0.0117567295209657 wvsat = -0.0835583479136885 pvsat = 9.09131850866372e-9   ua = -9.79958183545329e-10 lua = 7.06539746632345e-16 wua = 5.81237969530193e-15 pua = -4.94010647562068e-21   ub = 2.91296841672006e-18 lub = -8.74941832116534e-25 wub = -7.58481896246377e-24 pub = 6.05622094149507e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0374132654117264 lu0 = 6.45069071100329e-09 wu0 = 2.91159409148736e-08 pu0 = -3.21181715219691e-14   a0 = 1.57815040322507 la0 = 1.77759060843328e-08 wa0 = -2.28994671194983e-06 pa0 = -1.08723536657611e-13   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.187569564345236 lags = -5.14231324018407e-08 wags = -1.83020915659361e-08 pags = 2.44815449063109e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.861752645390261+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.02811969417008e-08 wnfactor = 2.94427209803226e-07 pnfactor = -3.64192284471693e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.149597251948763 lpclm = 1.05074756549794e-07 wpclm = -2.63897856427888e-06 ppclm = 4.86237165579067e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.82477577424507e-05 lalpha0 = -6.2392586619698e-11 walpha0 = -2.28205233045557e-10 palpha0 = 4.21491870561881e-16   alpha1 = 0.0   beta0 = 32.7088199111632 lbeta0 = -5.8010504044397e-06 wbeta0 = -4.08969951694548e-05 pbeta0 = 7.55361775200506e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 3508.266473688 lat = 0.0047598999914529 wat = 0.0397668978069747 pat = 5.39544125143218e-8   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.1226844289468e-18 lub1 = -1.16326054231727e-24 wub1 = -4.381820911013e-24 pub1 = 8.09316187714825e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.37 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.739664736334792+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.98791588951777e-08 wvth0 = 2.16085663906103e-07 pvth0 = -1.16753793884966e-13   k1 = 0.88325   k2 = -0.028041037072947 lk2 = 3.58209085470939e-09 wk2 = -1.86632756274018e-08 pk2 = 1.4633205166399e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 188420.07137475 lvsat = -0.0648136687382219 wvsat = -0.505830688445526 pvsat = 3.66750079126362e-7   ua = -1.32405787925235e-10 lua = -1.13252667243359e-17 wua = -1.23685313777182e-16 pua = 8.76574821591959e-23   ub = 1.3607074664663e-18 lub = 4.39801461095092e-25 wub = -3.95225900602975e-25 pub = -3.32637275981646e-32   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.044859423527802 lu0 = 1.4389903290078e-10 wu0 = -9.74944554778361e-09 pu0 = 8.00266696491525e-16   a0 = 3.14199757155161 la0 = -1.3067807516279e-06 wa0 = -1.02413817121257e-05 pa0 = 6.62603058840136e-12   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.0188307806233641 lags = 9.14962550676118e-08 wags = 1.14656916868022e-06 pags = -7.41814200167738e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.822003313839229+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.66140696086177e-08 wnfactor = 1.42646691677815e-07 pnfactor = 9.21367454778074e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -3.7727349440515 lpclm = 3.42723521391127e-06 wpclm = 2.43148430102153e-05 ppclm = -1.79671378643039e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -0.000140590561501121 lalpha0 = 9.75508260431375e-11 walpha0 = 9.79582670044057e-10 palpha0 = -6.01487574324379e-16   alpha1 = 0.0   beta0 = -5.26747557581609 lbeta0 = 2.63643402048949e-05 wbeta0 = 0.000204484975847273 pbeta0 = -1.32298916583524e-10   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.379199859999999 lkt1 = 5.47988084196013e-9   kt2 = -0.019151   at = -55156.2071053201 lat = 0.0544478878102426 wat = 0.4381820911013 pat = -2.83497678393265e-7   ute = -1.465198895 lute = 1.41106931680469e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -1.28362372552642e-17 lub1 = 7.063982711834e-24 wub1 = 1.13098426045092e-23 pub1 = -5.19745743720988e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.38 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.759172660767401+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.72578048982221e-08 wvth0 = 1.15253027314997e-07 pvth0 = -5.15164896674177e-14   k1 = 0.88325   k2 = -0.0139123907078416 lk2 = -5.55894554246468e-09 wk2 = 1.27916356066445e-08 pk2 = -5.71768203327165e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 55163.2823182108 lvsat = 0.0214016081863121 wvsat = 0.197423526658728 pvsat = -8.82455524870782e-8   ua = -3.02712926475661e-10 lua = 9.88610676178501e-17 wua = 3.81740786987641e-17 pua = -1.70632787412462e-23   ub = 1.3995151688713e-18 lub = 4.14693420946893e-25 wub = -1.44484676062839e-24 pub = 6.45826274146237e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0413898184832965 lu0 = 2.38868492222523e-09 wu0 = -2.75374404034359e-08 pu0 = 1.23088503361703e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.708250167194842+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.69826237262451e-08 wnfactor = 9.22135789698349e-07 pnfactor = -4.12181788094103e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.63860443699584 lpclm = -7.20811606875026e-07 wpclm = -1.11788742224835e-05 ppclm = 4.99680027321101e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -6.4930094011327e-06 lalpha0 = 1.07915872001747e-11 walpha0 = 1.61443495183728e-10 palpha0 = -7.21629821381938e-17   alpha1 = 0.0   beta0 = 32.1787734599999 lbeta0 = 2.13714132620842e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.65799999994 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -3.1939647150018e-18 lub1 = 8.25567370099795e-25 wub1 = 1.05992619505558e-23 pub1 = -4.73772170223111e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.39 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.93076736746378+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.94426266691647e-08 wvth0 = -2.96192657557197e-07 pvth0 = 1.32393971230865e-13   k1 = 0.88325   k2 = 0.00859077484697279 lk2 = -1.5617545501149e-08 wk2 = -8.05165333351456e-08 pk2 = 3.59897631693434e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 104476.749537704 lvsat = -0.000640821272260061 wvsat = -0.0539974173951911 pvsat = 2.41360896118067e-8   ua = 1.66630621568595e-10 lua = -1.1092892754826e-16 wua = -6.82487719912298e-17 pua = 3.05062455972718e-23   ub = -2.11537601382334e-19 lub = 1.13481145451148e-24 wub = 2.38450048558677e-24 pub = -1.06583833405049e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0333998941935409 lu0 = 5.96006922080595e-09 wu0 = 3.72006010511741e-08 pu0 = -1.66281478614601e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.2277700740348+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.8523550135252e-07 wnfactor = -1.86032923706131e-06 pnfactor = 8.31541124357086e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.128000232000002 lpclm = 4.01393324299249e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.869456438e-05 lalpha0 = -4.93676565395868e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.440127200000002 lkt1 = 3.10195768392001e-8   kt2 = -0.019151   at = 115413.814737024 lat = -0.0344240969940434 wat = -0.574434244959424 pat = 2.56764065417433e-7   ute = -1.30083493 lute = 7.75489420980013e-10   ua1 = -1.432830022e-09 lua1 = 1.53965669641369e-15   ub1 = 6.30577623000001e-18 lub1 = -3.42068383594278e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.40 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793874746824+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.72061228741093e-9   k1 = 0.88325   k2 = -0.042245136202 wk2 = 1.14570139832642e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 132965.844564 wvsat = -0.162479956463874   ua = 3.903402534698e-10 wua = -1.59195099345307e-15   ub = 1.192566965946e-18 wub = 1.72332402078016e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04544146501842 wu0 = -1.48965371255337e-8   a0 = 0.6263333686358 wa0 = 9.93177975511599e-7   keta = -0.012287877534 wketa = -5.33561131056816e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1077879014702 wags = 1.65431805172166e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.98447815154+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.82520568255446e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.821222460640001 wpclm = 5.08829227551036e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.14478230599999e-06 walpha0 = 2.75686689642077e-11   alpha1 = 0.0   beta0 = 21.60639121 wbeta0 = 6.48717682353732e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 208780.3136 wat = -0.281477502851789   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.41 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793874746824+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.72061228741009e-9   k1 = 0.88325   k2 = -0.042245136202 wk2 = 1.14570139832642e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 132965.844564 wvsat = -0.162479956463874   ua = 3.903402534698e-10 wua = -1.59195099345307e-15   ub = 1.192566965946e-18 wub = 1.72332402078017e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04544146501842 wu0 = -1.48965371255337e-8   a0 = 0.6263333686358 wa0 = 9.93177975511599e-7   keta = -0.012287877534 wketa = -5.33561131056815e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1077879014702 wags = 1.65431805172166e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.98447815154+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.82520568255446e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.82122246064 wpclm = 5.08829227551036e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.14478230599999e-06 walpha0 = 2.75686689642078e-11   alpha1 = 0.0   beta0 = 21.60639121 wbeta0 = 6.48717682353737e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 208780.3136 wat = -0.281477502851789   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.42 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.790910371669375+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.32614103370918e-08 wvth0 = 5.1224474484065e-09 pvth0 = -3.15319488263207e-15   k1 = 0.88325   k2 = -0.0437345759996019 lk2 = 1.16876132396251e-08 wk2 = 1.0983976451637e-08 pk2 = 3.71191888815319e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 138118.583119358 lvsat = -0.0404334673055531 wvsat = -0.200562650142707 pvsat = 2.98834364140097e-7   ua = 3.91171012000758e-10 lua = -6.51895056180834e-18 wua = -1.5945593971297e-15 pua = 2.04681071328815e-23   ub = 1.16541618945931e-18 lub = 2.13051762980167e-25 wub = 1.77329257553685e-24 pub = -3.92102549615882e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0447425074992988 lu0 = 5.48470986713865e-09 wu0 = -1.3066424708091e-08 pu0 = -1.43608665180989e-14   a0 = 0.628541395664266 la0 = -1.73263571799924e-08 wa0 = 9.93426126347864e-07 pa0 = -1.94723613805361e-15   keta = -0.012287877534 wketa = -5.33561131056816e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.101060657688965 lags = 5.27885877699355e-08 wags = 1.52148685692407e-07 pags = 1.04232452593997e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05049132061744+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.18004413566281e-07 wnfactor = -2.34119046039087e-08 pnfactor = 3.26936522041468e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.821222460640001 wpclm = 5.08829227551036e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -7.40231741073288e-06 lalpha0 = 9.84569158178068e-11 walpha0 = 6.6321087911366e-11 palpha0 = -3.04089688944485e-16   alpha1 = 0.0   beta0 = 16.919792259868 lbeta0 = 3.67756763493001e-05 wbeta0 = 1.20987695981303e-05 pbeta0 = -4.40340899399332e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414270958 lkt1 = 9.0561735852588e-8   kt2 = -0.019151   at = 304192.523289482 lat = -0.748698273662433 wat = -0.411192712716754 pat = 1.01787343579744e-6   ute = -1.33706986 lute = 3.01872452841962e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.43 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.802025951054856+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.95000679407443e-08 wvth0 = -4.46349603936867e-09 pvth0 = 3.37237955116176e-14   k1 = 0.88325   k2 = -0.04433723689548 lk2 = 1.40060412688157e-08 wk2 = 1.01556694846526e-08 pk2 = 6.89840419384426e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 145114.62716367 lvsat = -0.0673471507994073 wvsat = -0.213009462238378 pvsat = 3.46717076016769e-7   ua = 4.64929971962164e-10 lua = -2.90268636907897e-16 wua = -1.81051692737097e-15 pua = 8.51253702565642e-22   ub = 1.1578599726666e-18 lub = 2.42120423194712e-25 wub = 1.92513683412744e-24 pub = -9.76245286594306e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0461561968407622 lu0 = 4.62667621799507e-11 wu0 = -1.89917594936885e-08 pu0 = 8.43381344740794e-15   a0 = 0.177918923741793 la0 = 1.71621198359115e-06 wa0 = 1.87850683268371e-06 pa0 = -3.40684032228215e-12   keta = -0.040651119625867 lketa = 1.09112995242023e-07 wketa = 3.05227296385335e-08 pketa = -3.22680733733197e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.0254356709520466 lags = 3.43716852997047e-07 wags = 4.76427266893084e-07 pags = -1.14326270938487e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.956988350196316+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.58299795397814e-07 wnfactor = 5.778237557219e-08 pnfactor = 1.45832629239406e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.821222460640001 wpclm = 5.08829227551036e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.16299789545806e-05 lalpha0 = -1.3229921847405e-11 walpha0 = -2.44766961223455e-11 palpha0 = 4.52081150642265e-17   alpha1 = 0.0   beta0 = 24.0804539612766 lbeta0 = 9.22871103324548e-06 wbeta0 = -9.92565901215652e-07 pbeta0 = 6.32809444735423e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577635e-8   kt2 = -0.019151   at = 178637.92618422 lat = -0.265691496362848 wat = -0.214296226365803 pat = 2.60415409356143e-7   ute = -1.22166028 lute = -1.42106585683919e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.44 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.786287389175503+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.56883551055378e-09 wvth0 = 4.7122521270288e-09 pvth0 = 1.67763171087581e-14   k1 = 0.88325   k2 = -0.0468283046933552 lk2 = 1.86070086165421e-08 wk2 = 2.24298320110069e-08 pk2 = -1.57718021540568e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123220.156094145 lvsat = -0.0269083692565896 wvsat = -0.070878221052153 pvsat = 8.42026633831897e-8   ua = 6.97983662872098e-10 lua = -7.20715541266872e-16 wua = -2.50569484347796e-15 pua = 2.13523758112441e-21   ub = 8.1643827159928e-19 lub = 8.72721525162231e-25 wub = 2.80832669818462e-24 pub = -2.6074846008498e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0472776665684575 lu0 = -2.02507212429715e-09 wu0 = -1.97849338545987e-08 pu0 = 9.89879538756831e-15   a0 = 1.11100586904119 la0 = -7.18654115959784e-09 wa0 = 2.58326245162077e-08 pa0 = 1.50230027643049e-14   keta = 0.0430598171687215 lketa = -4.54999330644667e-08 wketa = -2.6630567940904e-07 pketa = 2.25557182179946e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.219173898878115 lags = -1.41149416472101e-08 wags = -1.74974511980456e-07 pags = 5.98672565696521e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.940233413235312+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.27353661399958e-07 wnfactor = -9.46261284811848e-08 pnfactor = 2.96079636191467e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.27853171664763 lpclm = 2.69162979351651e-06 wpclm = 9.39800459677578e-06 ppclm = -7.95997832140473e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.04693935335192e-05 lalpha0 = 4.60571697469005e-11 walpha0 = 6.28737707120187e-11 palpha0 = -1.16126974272308e-16   alpha1 = 0.0   beta0 = 21.5521891921279 lbeta0 = 1.38983806661562e-05 wbeta0 = 1.44098595470647e-05 pbeta0 = -2.21199697216632e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 31326.276947376 lat = 0.0063910574145138 wat = -0.0981355480583226 pat = 4.58682627717225e-8   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.0065958e-18 lub1 = 4.69311385258803e-25 wub1 = 5.87747175411144e-39   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.45 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.762307674893783+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.98793177911709e-08 wvth0 = 1.03837643444115e-07 pvth0 = -6.71815015813312e-14   k1 = 0.88325   k2 = -0.0350595707883207 lk2 = 8.63905576125245e-09 wk2 = 1.61297577080897e-08 pk2 = -1.04357274205261e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 62004.7466297314 lvsat = 0.0249402255440365 wvsat = 0.120849012235553 pvsat = -7.81876190302315e-8   ua = -1.70416530027428e-10 lua = 1.48072645163254e-17 wua = 6.47456421319527e-17 pua = -4.18895240203832e-23   ub = 1.51182378195509e-18 lub = 2.83739733288006e-25 wub = -1.14435602030604e-24 pub = 7.40382324153725e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.049810575936172 lu0 = -4.17041089802012e-09 wu0 = -3.42938329910145e-08 pu0 = 2.21876298315246e-14   a0 = 1.03886093318061 la0 = 5.39192094852069e-08 wa0 = 1.8451437036396e-07 pa0 = -1.19378214424296e-13   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.339213878839846 lags = -1.15787124115076e-07 wags = -4.4166852717313e-07 pags = 2.85753353721635e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.632986117612829+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.32880496530146e-07 wnfactor = 1.07966315066851e-06 pnfactor = -6.98526943198419e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.1321132135 lpclm = -1.97138713289512e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 0.000120428427757596 lalpha0 = -6.48114523171761e-11 walpha0 = -3.14368853560094e-10 palpha0 = 2.03392247089431e-16   alpha1 = 0.0   beta0 = 45.9821296461993 lbeta0 = -6.79343687927597e-06 wbeta0 = -4.95751021166654e-05 pbeta0 = 3.20743970180529e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37919986 lkt1 = 5.47988084196013e-9   kt2 = -0.019151   at = 70806.9071053201 lat = -0.0270484836004426 wat = -0.18625586268002 pat = 1.20504935571895e-7   ute = -1.465198895 lute = 1.41106931680469e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -1.0554788815e-17 lub1 = 6.01553919426159e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.46 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.792920770841267+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.00730732964922e-08 wvth0 = -5.20467487390611e-08 pvth0 = 3.36735177796929e-14   k1 = 0.88325   k2 = -0.0058062623341657 lk2 = -1.02874252622675e-08 wk2 = -2.73929394292063e-08 pk2 = 1.77228483095444e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 91765.2953348487 lvsat = 0.00568556717950763 wvsat = 0.0159760747152458 pvsat = -1.03362966757179e-8   ua = -5.10383846218894e-10 lua = 2.34761358549777e-16 wua = 1.06766279050925e-15 pua = -6.90762878180416e-22   ub = 1.28756789446683e-18 lub = 4.28830152910481e-25 wub = -8.89889641644923e-25 pub = 5.75746139689285e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03089042582787 lu0 = 8.07066133994969e-09 wu0 = 2.45112828024508e-08 pu0 = -1.58584568152265e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.975593975513654+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.87819910216772e-08 wnfactor = -4.03169810030958e-07 pnfactor = 2.60845222712689e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.23882855337614 lpclm = -2.66182044174613e-07 wpclm = -4.23975403640844e-06 ppclm = 2.74306150499975e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.79838674904791e-05 lalpha0 = -5.00111604819516e-12 walpha0 = -9.46900244607457e-12 palpha0 = 6.12631201657597e-18   alpha1 = 0.0   beta0 = 32.17877346 lbeta0 = 2.13714132620845e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -1.60443453858052e-18 lub1 = 2.24785282378057e-25 wub1 = 2.71947129074112e-24 pub1 = -1.75945985251143e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.47 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.876998027230725+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.75082832280058e-08 wvth0 = -2.96414770651607e-08 pvth0 = 2.36586750152608e-14   k1 = 0.88325   k2 = -0.0114940857020103 lk2 = -7.74504784636807e-09 wk2 = 1.90503065432129e-08 pk2 = -3.03663243468337e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110240.376059935 lvsat = -0.00257253525347589 wvsat = -0.0825694892628603 pvsat = 3.37121907845996e-8   ua = 5.95321779863884e-10 lua = -2.59473576430459e-16 wua = -2.19340288053773e-15 pua = 7.66887821858189e-22   ub = -6.2489136925669e-19 lub = 1.28367266936521e-24 wub = 4.43362242590048e-24 pub = -1.80378922533456e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0438080717040657 lu0 = 2.29665448033251e-09 wu0 = -1.43959405871703e-08 pu0 = 1.53252733880667e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.03657748603187+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.16040766454171e-07 wnfactor = -9.12528691013654e-07 pnfactor = 4.88521511487622e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.58250637215227 lpclm = 9.94915168847628e-07 wpclm = 8.4795080728169e-06 ppclm = -2.94227058815444e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.48743448390417e-05 lalpha0 = -3.61120295631972e-12 walpha0 = 1.8938004892149e-11 palpha0 = -6.57122256550721e-18   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768392001e-8   kt2 = -0.019151   at = -462.432000000088 lat = 0.017370963029952   ute = -1.30083493 lute = 7.75489420980013e-10   ua1 = -1.432830022e-09 lua1 = 1.53965669641369e-15   ub1 = 7.40293270716105e-18 lub1 = -3.80138177332698e-24 wub1 = -5.43894258148224e-24 pub1 = 1.8872369305782e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.48 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.788888825533334+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.94655172076689e-8   k1 = 0.88325   k2 = -0.041005812864 wk2 = 7.7919531612101e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 40953.9706346667 wvsat = 0.109627494402335   ua = -1.47719457254667e-10 wua = -7.42706449916182e-19   ub = 1.78259239769333e-18 wub = -2.15629087296765e-26   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0416061119076 wu0 = -3.55421668808073e-9   a0 = 0.809344787270934 wa0 = 4.51956843090571e-7   keta = -0.0350448771493333 wketa = 1.39433439127407e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.158104925658933 wags = 1.66288670026311e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.996488947386667+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.72675658181688e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.34623864050667 wpclm = -1.32155777859949e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 20.9825378666667 wbeta0 = 8.33210330660372e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414388464 wkt1 = 3.4477668854912e-8   kt2 = -0.019151   at = 155959.085866667 wat = -0.12526886350618   ute = -1.410812716 wute = 3.31847562728527e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.49 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.788888825533333+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.94655172076689e-8   k1 = 0.88325   k2 = -0.041005812864 wk2 = 7.79195316121013e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 40953.9706346667 wvsat = 0.109627494402335   ua = -1.47719457254667e-10 wua = -7.4270644991628e-19   ub = 1.78259239769333e-18 wub = -2.15629087296765e-26   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0416061119076 wu0 = -3.55421668808075e-9   a0 = 0.809344787270934 wa0 = 4.51956843090571e-7   keta = -0.0350448771493333 wketa = 1.39433439127407e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.158104925658933 wags = 1.66288670026311e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.996488947386667+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.72675658181684e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.34623864050667 wpclm = -1.32155777859949e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 20.9825378666667 wbeta0 = 8.33210330660375e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414388464 wkt1 = 3.44776688549118e-8   kt2 = -0.019151   at = 155959.085866667 wat = -0.12526886350618   ute = -1.410812716 wute = 3.31847562728527e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.50 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.783312335400814+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.37586399990177e-08 wvth0 = 2.75921808897094e-08 pvth0 = -6.37698161396889e-14   k1 = 0.88325   k2 = -0.0442576593710625 lk2 = 2.55171940150683e-08 wk2 = 1.25308950907243e-08 pk2 = -3.71864109757111e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 25724.331483223 lvsat = 0.119506765206431 wvsat = 0.131821769374847 pvsat = -1.74158164989453e-7   ua = -1.47820520472641e-10 lua = 7.93041656561362e-19 wua = -5.95426213856153e-19 pua = -1.15570595043995e-24   ub = 1.76237596185759e-18 lub = 1.58638088972977e-25 wub = 7.89866494523938e-27 pub = -2.31184556165031e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.041448165077257 lu0 = 1.23940656644618e-09 wu0 = -3.3240395086472e-09 pu0 = -1.80619710453454e-15   a0 = 0.81386343182544 la0 = -3.54577405581959e-08 wa0 = 4.4537178623213e-07 pa0 = 5.16728489773854e-14   keta = -0.0350448771493333 wketa = 1.39433439127407e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.13598649143763 lags = 1.73563043676485e-07 wags = 4.88622381408097e-08 pags = -2.52934812054092e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.09886048844574+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.03308049488942e-07 wnfactor = -1.66454431575879e-07 pnfactor = 1.17066724698463e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.34623864050667 wpclm = -1.32155777859949e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.55648537187109e-05 lalpha0 = -8.61484276077233e-12 walpha0 = -1.59991100710713e-12 palpha0 = 1.25544792740156e-17   alpha1 = 0.0   beta0 = 15.4837886710508 lbeta0 = 4.3148607955509e-05 wbeta0 = 1.63454744993683e-05 pbeta0 = -6.28808115624268e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.437141908947376 lkt1 = 1.78545963953829e-07 wkt1 = 6.76364462042822e-08 pkt1 = -2.60196461637628e-13   kt2 = -0.019151   at = 257591.139964946 lat = -0.797505305660442 wat = -0.273378069000036 pat = 1.16221086198141e-6   ute = -1.48665753249125 lute = 5.95153213179435e-07 wute = 4.42376820559764e-07 pute = -8.67321538792096e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.51 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.799451986452162+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.83303716404023e-08 wvth0 = 3.14851007189787e-09 pvth0 = 3.02646432850429e-14   k1 = 0.88325   k2 = -0.0426496486975625 lk2 = 1.93311994662632e-08 wk2 = 5.16495140624559e-09 pk2 = -8.84972874473287e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 26688.5218524671 lvsat = 0.115797538354613 wvsat = 0.137213006407287 pvsat = -1.9489817837593e-7   ua = -1.46539998021917e-10 lua = -4.13311028406069e-18 wua = -2.21189337729186e-18 pua = 5.06282059675614e-24   ub = 1.83196617111776e-18 lub = -1.09074471787974e-25 wub = -6.84028194017736e-26 pub = 6.23461858971499e-32   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0411916969960788 lu0 = 2.22603568418526e-09 wu0 = -4.31020438700775e-09 pu0 = 1.98756537621032e-15   a0 = 0.511662757202588 la0 = 1.12710402390647e-06 wa0 = 8.91523524039429e-07 pa0 = -1.66466664024296e-12   keta = -0.0272983732800593 lketa = -2.98006919340432e-08 wketa = -8.96545395189446e-09 pketa = 8.81298246620812e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.209181391132396 lags = -1.08016710720681e-07 wags = -6.69654213620244e-08 pags = 1.92652572466079e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.938436254583346+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.86158267759599e-07 wnfactor = 1.12646636345191e-07 pnfactor = 9.69693461072252e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.34623864050667 wpclm = -1.32155777859949e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.12332215668925e-05 lalpha0 = 8.04888548442276e-12 walpha0 = 6.26971767432347e-12 palpha0 = -1.77198720886464e-17   alpha1 = 0.0   beta0 = 22.7839113918934 lbeta0 = 1.50651380501456e-05 wbeta0 = 2.84170981156178e-06 pbeta0 = -1.09320178611407e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.3947963557764e-8   kt2 = -0.019151   at = 96459.2633333333 lat = -0.1776332321049 wat = 0.0287313907124267   ute = -1.26953070924909 lute = -2.40130636057655e-07 wute = 1.41567603381759e-07 pute = 2.8988730836265e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.52 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.780343001364874+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.69636562900265e-08 wvth0 = 2.22916377545046e-08 pvth0 = -5.09244554094127e-15   k1 = 0.88325   k2 = -0.0387719097183175 lk2 = 1.21690698599434e-08 wk2 = -1.39540929983206e-09 pk2 = 3.26716563434259e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 81147.4832575212 lvsat = 0.0152125990649383 wvsat = 0.0535436309089786 pvsat = -4.03620132018112e-8   ua = -1.49607582925674e-10 lua = 1.53267608699014e-18 wua = 8.93528449761271e-19 pua = -6.72850041905429e-25   ub = 1.75526190927161e-18 lub = 3.25972259821927e-26 wub = 3.19360439071176e-26 pub = -1.22978289890285e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419217928954986 lu0 = 8.77558779299509e-10 wu0 = -3.94596579456816e-09 pu0 = 1.31482179531473e-15   a0 = 1.12748943513215 la0 = -1.03192286559339e-08 wa0 = -2.29143573531125e-08 pa0 = 2.42873245587211e-14   keta = -0.0711915344450867 lketa = 5.12693622335062e-08 wketa = 7.15707567292875e-08 pketa = -6.06194289591123e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.128832671522715 lags = 4.03862495163244e-08 wags = 9.21923224074878e-08 pags = -1.01309552067798e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.862817868854418+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.64921679756705e-08 wnfactor = 1.34315480240787e-07 pnfactor = 5.69472947958753e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.93616928976111 lpclm = -1.08959365014387e-06 wpclm = -3.06616440708485e-06 ppclm = 3.22226401831966e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.02484532040256e-05 lalpha0 = -8.60212113611905e-12 walpha0 = -2.79683631876964e-11 palpha0 = 4.55173839303722e-17   alpha1 = 0.0   beta0 = 29.5636774592696 lbeta0 = 2.54300504042671e-06 wbeta0 = -9.28257879725952e-06 pbeta0 = 1.14613734593116e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = -19801.98715792 lat = 0.037099669894938 wat = 0.0530664764063821 pat = -4.4946562585536e-8   ute = -1.48504006301079 lute = 1.57912123209256e-07 wute = 5.5136068986231e-07 pute = -4.66994785263718e-13   ua1 = 3.0044e-9   ub1 = -4.2534596947376e-18 lub1 = 9.2526554274462e-25 wub1 = 7.30052570818664e-25 pub1 = -1.34839687756608e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.53 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.802984306331764+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.21321203866009e-09 wvth0 = -1.64556841204789e-08 pvth0 = 2.77259936246626e-14   k1 = 0.88325   k2 = -0.0251924467891824 lk2 = 6.67454871446972e-10 wk2 = -1.30503670315539e-08 pk2 = 1.31387516637028e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 116468.503797368 lvsat = -0.0147038108380241 wvsat = -0.040217092546355 pvsat = 3.90520069147275e-8   ua = -1.37880000893315e-10 lua = -8.40042170826954e-18 wua = -3.14748957685915e-17 pua = 2.67427521131004e-23   ub = 8.33320036528148e-19 lub = 8.1346908500969e-25 wub = 8.62188534075005e-25 pub = -8.26190525527626e-31   uc = 6.49562847471529e-11 luc = 1.05679735114796e-18 wuc = 3.6898782989667e-18 puc = -3.12527526092865e-24   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0360892389134166 lu0 = 5.81765034636724e-09 wu0 = 6.28438675707609e-09 pu0 = -7.35014359099224e-15   a0 = 1.09300424424452 la0 = 1.88892452332168e-08 wa0 = 2.43959234081893e-08 pa0 = -1.57838209021718e-14   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.229131060693314 lags = -4.45650819337243e-08 wags = -1.16119728405847e-07 pags = 7.51278386023854e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.19404169184913+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.27034108918671e-07 wnfactor = -5.79550987465098e-07 pnfactor = 6.61582198812212e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.70475735929648 lpclm = -4.66049848073503e-08 wpclm = 1.26382288648291e-06 ppclm = -4.45174599510122e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.54370765068824e-05 lalpha0 = -4.52695243291255e-12 walpha0 = -3.87709057554809e-12 palpha0 = 2.51124133056992e-17   alpha1 = 0.0   beta0 = 27.778489982421 lbeta0 = 4.05503384069277e-06 wbeta0 = 4.25866709014364e-06 pbeta0 = -7.8722298763821e-15   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37919986 lkt1 = 5.47988084196013e-9   kt2 = -0.019151   at = 7825.35000000001 lat = 0.0136997021049   ute = -1.465198895 lute = 1.41106931680469e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -1.1030813524182e-17 lub1 = 6.66558935333044e-24 wub1 = 1.4077516806617e-24 pub1 = -1.92239853581559e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.54 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.762223799128151+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.41582654749769e-08 wvth0 = 3.8733651283908e-08 pvth0 = -7.98073373127966e-15   k1 = 0.88325   k2 = -0.0125117238921877 lk2 = -7.53679531278807e-09 wk2 = -7.5628243199754e-09 pk2 = 9.58838835490944e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 78561.0039800616 lvsat = 0.00982181083877542 wvsat = 0.0550252311730881 pvsat = -2.25684431392198e-8   ua = -1.54523843871962e-10 lua = 2.3679116851131e-18 wua = 1.52751586886452e-17 pua = -3.50387861996937e-24   ub = 9.83392559704077e-19 lub = 7.16374263530187e-25 wub = 9.65050925163861e-27 pub = -2.74610358999256e-31   uc = 5.25021707717075e-11 luc = 9.11443473566546e-18 wuc = 4.05205291914631e-17 puc = -2.69541907592613e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0424830326312896 lu0 = 1.68095532401546e-09 wu0 = -9.77162603815612e-09 pu0 = 3.03787190334382e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.702012659859722+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.69821362797095e-09 wnfactor = 4.0589440340294e-07 pnfactor = 2.40128271560625e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.179613658207871 lpclm = 2.93155637785162e-07 wpclm = -1.10732935320818e-06 ppclm = 1.08892770343866e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.02933029400651e-05 lalpha0 = 1.21202428439503e-11 walpha0 = 1.03728379885537e-10 palpha0 = -4.45068196060368e-17   alpha1 = 0.0   beta0 = 27.5336270022971 lbeta0 = 4.21345676075122e-06 wbeta0 = 1.37371287805364e-05 pbeta0 = -6.14030424509686e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.65800000002 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = 3.99711575947093e-19 lub1 = -7.29800359101699e-25 wub1 = -3.20740604692031e-24 pub1 = 1.06354390172178e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.55 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.860278806730389+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.96709501531172e-08 wvth0 = 1.9802407474242e-08 pvth0 = 4.81267214227858e-16   k1 = 0.88325   k2 = -0.0130754449860965 lk2 = -7.28481987590616e-09 wk2 = 2.37268730049153e-08 pk2 = -4.39766829355417e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 86583.0210305767 lvsat = 0.00623608152543387 wvsat = -0.0126074039756978 pvsat = 7.66239791539551e-9   ua = -1.52594375186884e-10 lua = 1.50546619544497e-18 wua = 1.84155481231457e-17 pua = -4.90758873173895e-24   ub = 1.0726955610575e-18 lub = 6.7645707216723e-25 wub = -5.8666498381313e-25 pub = -8.06568201620602e-33   uc = 9.61030889622792e-11 luc = -1.03745652826654e-17 wuc = -8.842081498086e-17 puc = 3.06807849069487e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0384543125386977 lu0 = 3.48173680332279e-09 wu0 = 1.43677422264578e-09 pu0 = -1.97212609563094e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.497451206703296+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.27378920726075e-08 wnfactor = 6.81833767854961e-07 pnfactor = -9.93282056028892e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.723671843871333 lpclm = 6.96911611217538e-07 wpclm = 5.93966985165545e-06 ppclm = -2.06098228314652e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.49943407398231e-05 lalpha0 = -3.65283985394826e-12 walpha0 = 1.8583140054801e-11 palpha0 = -6.44808943505516e-18   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768391999e-8   kt2 = -0.019151   at = -462.43200000003 lat = 0.017370963029952   ute = -1.30083493 lute = 7.75489420979166e-10   ua1 = -1.43283002200001e-09 lua1 = 1.53965669641369e-15   ub1 = 6.14110821226189e-18 lub1 = -3.2961242759815e-24 wub1 = -1.70733890812099e-24 pub1 = 3.93034891618429e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.56 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7976509216+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.69644451294716e-9   k1 = 0.88325   k2 = -0.033177657664 wk2 = -3.61608003699151e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 124374.55648 wvsat = -0.0119419927147558   ua = -1.477422131512e-10 wua = -7.09544099851084e-19   ub = 1.738915932256e-18 wub = 4.20871537638739e-26   uc = 9.2162363728e-11 wuc = -3.78293311277242e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04034103277728 wu0 = -1.71060675083235e-9   a0 = 1.11509733491568 wa0 = 6.38120938750018e-9   keta = -0.032444287624 wketa = 1.01534839927562e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1897184365704 wags = -2.94417553567364e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.794767531280001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.76702667645406e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.68718920056 wpclm = 1.64177288160969e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.6833142368e-05 walpha0 = 4.56139478740254e-11   alpha1 = 0.0   beta0 = 26.190712144 wbeta0 = 7.42189266851649e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.386900768 wkt1 = -5.58037042745575e-9   kt2 = -0.019151   at = -83169.28 wat = 0.22321481709824   ute = -1.2106704704 wute = 4.01786670776829e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.57 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7976509216+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.69644451294716e-9   k1 = 0.88325   k2 = -0.033177657664 wk2 = -3.61608003699151e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 124374.55648 wvsat = -0.0119419927147558   ua = -1.477422131512e-10 wua = -7.09544099851084e-19   ub = 1.738915932256e-18 wub = 4.20871537638739e-26   uc = 9.2162363728e-11 wuc = -3.78293311277242e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04034103277728 wu0 = -1.71060675083235e-9   a0 = 1.11509733491568 wa0 = 6.38120938749934e-9   keta = -0.032444287624 wketa = 1.01534839927562e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1897184365704 wags = -2.94417553567364e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.79476753128+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.76702667645406e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.687189200560001 wpclm = 1.64177288160969e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.6833142368e-05 walpha0 = 4.56139478740254e-11   alpha1 = 0.0   beta0 = 26.190712144 wbeta0 = 7.42189266851649e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.386900768 wkt1 = -5.58037042745618e-9   kt2 = -0.019151   at = -83169.2800000001 wat = 0.22321481709824   ute = -1.2106704704 wute = 4.01786670776829e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.58 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.800700238992214+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.39279508862563e-08 wvth0 = 2.25264988273585e-09 pvth0 = 3.48703942501473e-14   k1 = 0.88325   k2 = -0.0295205023061041 lk2 = -2.8697646893234e-08 wk2 = -8.94568179729601e-09 pk2 = 4.1821310398685e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 124374.55648 wvsat = -0.0119419927147558   ua = -1.45758867883595e-10 lua = -1.55632825480606e-17 wua = -3.59988902509347e-18 pua = 2.26804961635488e-23   ub = 1.81457804073792e-18 lub = -5.93719505988109e-25 wub = -6.81758422236983e-26 pub = 8.65232185832515e-31   uc = 9.2162363728e-11 wuc = -3.78293311277242e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.040769927738821 lu0 = -3.36553275868228e-09 wu0 = -2.33563880944566e-09 pu0 = 4.90461781348973e-15   a0 = 1.10970722449489 la0 = 4.22961210104272e-08 wa0 = 1.42362604246071e-08 pa0 = -6.16384755174637e-14   keta = -0.032444287624 wketa = 1.01534839927562e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.209586691238423 lags = -1.55905916224412e-07 wags = -5.83959218304837e-08 pags = 2.27202938961165e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.670272151516978+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.76913502065122e-07 wnfactor = 4.58130780537098e-07 pnfactor = -1.42366386186752e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.68718920056 wpclm = 1.64177288160969e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -3.36154362765962e-05 lalpha0 = 1.3169042534864e-10 walpha0 = 7.00709190453739e-11 palpha0 = -1.91913510383976e-16   alpha1 = 0.0   beta0 = 28.2604179102127 lbeta0 = -1.624095217159e-05 wbeta0 = -2.27400950389618e-06 pbeta0 = 2.36680695272754e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.383218017526312 lkt1 = -2.88984914085244e-08 wkt1 = -1.09472721547649e-08 pkt1 = 4.21140027175722e-14   kt2 = -0.019151   at = -285720.55605284 lat = 1.58941702746877 wat = 0.518394412100252 pat = -2.31627014946646e-6   ute = -1.2106704704 wute = 4.01786670776838e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.59 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.790209748693623+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.64288184255533e-08 wvth0 = 1.6617297095317e-08 pvth0 = -2.03902024715924e-14   k1 = 0.88325   k2 = -0.0404658281494685 lk2 = 1.34088683916272e-08 wk2 = 1.98245225094388e-09 pk2 = -2.19068291017239e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 134607.819722117 lvsat = -0.0393672204267395 wvsat = -0.0200586497325369 pvsat = 3.12246659142059e-8   ua = -1.48757911528824e-10 lua = -4.02600363147475e-18 wua = 1.02028971963273e-18 pua = 4.90673321508917e-24   ub = 1.58737260741686e-18 lub = 2.80336615121946e-25 wub = 2.88045337728062e-25 pub = -5.05145706345376e-31   uc = 1.15432781536208e-10 luc = -8.95209715223262e-17 wuc = -7.17414971629679e-17 puc = 1.30459627967258e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0397551260167555 lu0 = 5.38395258879452e-10 wu0 = -2.21667800627198e-09 pu0 = 4.44697726913188e-15   a0 = 1.13201101245189 la0 = -4.35062390071515e-08 wa0 = -1.25149511214264e-08 pa0 = 4.12730607831689e-14   keta = -0.0556837992318222 lketa = 8.94020758021295e-08 wketa = 3.24008543710173e-08 pketa = -8.55853223819851e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.13707813714414 lags = 1.2303347625654e-07 wags = 3.81112275010932e-08 pags = -1.44058713417321e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.972141368539509+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.8437314965152e-07 wnfactor = 6.35279041359614e-08 pnfactor = 9.43678792073784e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.687189200560001 wpclm = 1.64177288160969e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -8.03605407933667e-06 lalpha0 = 3.3286900147133e-11 walpha0 = 3.43509872277784e-11 palpha0 = -5.44994327607313e-17   alpha1 = 0.0   beta0 = 20.9215116206291 lbeta0 = 1.19917175797499e-05 wbeta0 = 5.55579989742336e-06 pbeta0 = -6.45309762226925e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.39479635577635e-8   kt2 = -0.019151   at = 226657.16421064 lat = -0.381692889096754 wat = -0.16100705181928 pat = 2.97377770611484e-7   ute = -1.17944759170522 lute = -1.20113977218519e-07 wute = 1.02887555201389e-08 pute = 1.14986071303107e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.60 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7907304906401+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.54670153407995e-08 wvth0 = 7.1538665338034e-09 pvth0 = -2.91137871250495e-15   k1 = 0.88325   k2 = -0.041801873307151 lk2 = 1.58765250932345e-08 wk2 = 3.02018087788382e-09 pk2 = -2.13573853677456e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 129101.287806358 lvsat = -0.0291967330697793 wvsat = -0.0163398320904778 pvsat = 2.43560617927695e-8   ua = -1.5584808691025e-10 lua = 9.06945103556243e-18 wua = 9.98786483051538e-18 pua = -1.16562524686593e-23   ub = 1.74451631587589e-18 lub = -9.90561438997265e-27 wub = 4.75956831274481e-26 pub = -6.10385605932045e-32   uc = 3.54002495842735e-11 luc = 5.82979945374493e-17 wuc = 4.48905519108415e-17 puc = -8.49581338233811e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0392238305150842 lu0 = 1.51969061232927e-09 wu0 = -1.42036338911726e-11 pu0 = 3.79037937985717e-16   a0 = 1.0924620965587 la0 = 2.95400549627539e-08 wa0 = 2.81312633686823e-08 pa0 = -3.37999283330622e-14   keta = -0.00441625104585688 lketa = -5.28836795167387e-09 wketa = -2.57413979706773e-08 pketa = 2.18026037015921e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.250695725391704 lags = -8.68166185904764e-08 wags = -8.53996809002204e-08 pags = 8.40642052471876e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.867688878150487+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.54913776214061e-09 wnfactor = 1.27216919425553e-07 pnfactor = -2.32648403862836e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.45698114832333 lpclm = 3.2687809504316e-06 wpclm = 3.33600887153911e-06 ppclm = -3.12923015409577e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -3.20605689453068e-06 lalpha0 = 2.43659629667569e-11 walpha0 = 6.21208201501044e-12 palpha0 = -2.52726877742178e-18   alpha1 = 0.0   beta0 = 20.5806993898891 lbeta0 = 1.26211929985554e-05 wbeta0 = 3.8083870070732e-06 pbeta0 = -3.22565047757289e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16612.056 lat = 0.00625748513678401   ute = -0.861661664767044 lute = -7.07060135270355e-07 wute = -3.57093636925486e-07 pute = 7.93536206796685e-13   ua1 = 3.0044e-9   ub1 = -3.02226967779659e-18 lub1 = -1.34872518188519e-24 wub1 = -1.06417049038961e-24 pub1 = 1.96550799736275e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.61 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.780892260890475+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.37998582035147e-08 wvth0 = 1.57392304374755e-08 pvth0 = -1.018306174382e-14   k1 = 0.88325   k2 = -0.0355965130214804 lk2 = 1.06206718063155e-08 wk2 = 2.11156192130382e-09 pk2 = -1.3661510012167e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 52789.8878868839 lvsat = 0.0354379543024166 wvsat = 0.0525822638489204 pvsat = -3.40199885585576e-8   ua = -1.48510246409012e-10 lua = 2.85440286078083e-18 wua = -1.59833539366026e-17 pua = 1.03410062300267e-23   ub = 1.49606048034243e-18 lub = 2.00532999925169e-25 wub = -1.03628416619107e-25 pub = 6.70461347547319e-32   uc = 2.28526513149174e-10 luc = -1.05277246934331e-16 wuc = -2.34682324113125e-16 puc = 1.51836178148655e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.039142367327192 lu0 = 1.58868879198937e-09 wu0 = 1.83503829465383e-09 pu0 = -1.18724408610492e-15   a0 = 1.14396233539311 la0 = -1.40799263266437e-08 wa0 = -4.98657104873773e-08 pa0 = 3.22624165653866e-14   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.109198222880707 lags = 3.30297850713033e-08 wags = 5.86593556011677e-08 pags = -3.79517818429769e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.50648522875654+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.14483571947721e-07 wnfactor = 4.22430546651439e-07 pnfactor = -2.73306649655828e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.61390052368908 lpclm = -1.0261848334195e-06 wpclm = -1.51838672013175e-06 ppclm = 9.82374950511158e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.39536728942978e-06 lalpha0 = 1.87746491028809e-11 walpha0 = 1.36713886007194e-11 palpha0 = -8.84519702522499e-18   alpha1 = 0.0   beta0 = 30.7007734600001 lbeta0 = 4.04963194220847e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37919986 lkt1 = 5.4798808419597e-9   kt2 = -0.019151   at = 7825.35000000003 lat = 0.0136997021049   ute = -3.15009630732366 lute = 1.23121196889011e-06 wute = 2.45541447815858e-06 pute = -1.58861879156591e-12   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -1.37159705200171e-17 lub1 = 7.70868971966376e-24 wub1 = 5.32085245194806e-24 pub1 = -3.44251704447607e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.62 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.788802704399999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.86819119990614e-8   k1 = 0.88325   k2 = -0.0177013092921 lk2 = -9.57274473741399e-10   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 116319.138275 lvsat = -0.00566458128918917   ua = -1.44042079764e-10 lua = -3.64384042086863e-20   ub = 9.900147077e-19 lub = 5.27937530184008e-25   uc = 8.03072258399999e-11 luc = -9.38144311531821e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0357777746911999 lu0 = 3.7655331231793e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.980536076599998+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.7793101048727e-9   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.580232134999999 lpclm = 1.04037427889511e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 6.088477327e-05 lalpha0 = -1.84201917148642e-11   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.65799999994 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.63 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.859982344799839+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.3134390744702e-08 wvth0 = 2.0234443817324e-08 pvth0 = -9.04451310413095e-15   k1 = 0.88325   k2 = 0.0235275055354845 lk2 = -1.93859774982641e-08 wk2 = -2.96148996137889e-08 pk2 = 1.3237445518769e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 96358.1329724207 lvsat = 0.00325770862698954 wvsat = -0.0268527528094429 pvsat = 1.20028045672816e-8   ua = -1.01298124906295e-10 lua = -1.91423878102345e-17 wua = -5.63388877807578e-17 pua = 2.51826940935698e-23   ub = -3.61931914548622e-19 lub = 1.13223874307643e-24 wub = 1.50402911340747e-24 pub = -6.72279957285548e-31   uc = -9.65165360983478e-11 luc = 6.9656302938456e-17 wuc = 1.92285305576992e-16 puc = -8.59488395986373e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.038996373468258 lu0 = 2.32686453021719e-09 wu0 = 6.46824493509839e-10 pu0 = -2.89121493055981e-16   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.23750544093995+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.07082398183983e-07 wnfactor = -3.96653188131988e-07 pnfactor = 1.77298421950364e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.35211025 lpclm = -7.17327714406501e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.774603088e-05 lalpha0 = -8.0774978089277e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768392003e-8   kt2 = -0.019151   at = -58287.0162196074 lat = 0.0432177426319374 wat = 0.0842682291799074 pat = -3.766671868821e-8   ute = -0.265785501988187 lute = -4.61877114208307e-07 wute = -1.50838581183703e-06 pute = 6.74227340489789e-13   ua1 = -1.43283002200001e-09 lua1 = 1.53965669641369e-15   ub1 = 1.82105969641511e-17 lub1 = -8.94499307781804e-24 wub1 = -1.92963014221591e-23 pub1 = 8.62517658748523e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.64 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7743732176+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.89803767737794e-8   k1 = 0.88325   k2 = -0.038262105184 wk2 = 1.25130224948469e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 142738.6288 wvsat = -0.0295220660592704   ua = -1.552993028112e-10 wua = 6.52491828838429e-18   ub = 1.5408392024e-18 wub = 2.3170759186886e-25   uc = 4.0321865408e-11 wuc = 1.17979926379984e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0376285567512 wu0 = 8.86068248742244e-10   a0 = 2.00952836416384 wa0 = -8.49864770359997e-7   keta = -0.026319503488 wketa = 4.29017914109029e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.1553244588784 wags = 3.48387463963672e-9   b0 = 1.52898095264e-07 wb0 = -1.14843545416989e-13   b1 = -9.68050021119999e-10 wb1 = 9.26722029618344e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.12537141808+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -3.97870780193284e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.35407942736 wpclm = -2.22696590604715e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.8592558768e-05 walpha0 = -7.44551922907654e-12   alpha1 = 0.0   beta0 = 21.98655168 wbeta0 = 4.76686571232254e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.398388464 wkt1 = 5.41689285491168e-9   kt2 = -0.019151   at = 404630.88 wat = -0.24376017847104   ute = -1.270552352 wute = 9.75040713884158e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.65 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.754577375960513+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.92887791877122e-07 wvth0 = 4.79310943419933e-08 pvth0 = -3.76114626266302e-13   k1 = 0.88325   k2 = -0.039116841523948 lk2 = 1.69639401726383e-08 wk2 = 2.0695481856076e-09 pk2 = -1.62397156387881e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 162904.486171066 lvsat = -0.400231488921552 wvsat = -0.0488270026474512 pvsat = 3.83144806196513e-7   ua = -1.59756327305937e-10 lua = 8.84585027487079e-17 wua = 1.07916634933922e-17 pua = -8.46820323493598e-23   ub = 1.382564973217e-18 lub = 3.14126641075585e-24 wub = 3.83224777659582e-25 pub = -3.00715946514786e-30   uc = 3.2262922774205e-11 luc = 1.59945721627732e-16 wuc = 1.95128828928713e-17 puc = -1.53117318880001e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0370233035182693 lu0 = 1.20124524404295e-08 wu0 = 1.46548201065263e-09 pu0 = -1.1499616820843e-14   a0 = 2.59005181768386 la0 = -1.15216408546835e-05 wa0 = -1.40560451660234e-06 pa0 = 1.10297589633153e-11   keta = -0.0292500280821072 lketa = 5.81620805919024e-08 wketa = 7.09559377922594e-09 pketa = -5.56790250472731e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.152944702700748 lags = 4.72309875412651e-08 wags = 5.76203426655188e-09 pags = -4.5214602221153e-14   b0 = 2.31345130516106e-07 lb0 = -1.55693721039006e-12 wb0 = -1.89941519840113e-13 pb0 = 1.49046844700409e-18   b1 = -1.60107293470569e-09 lb1 = 1.25635969036145e-14 wb1 = 1.53271992897724e-15 pb1 = -1.20272318246054e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.15254907356449+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.39394547913535e-07 wnfactor = -6.58044650358768e-08 pnfactor = 5.16366715874011e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 4.87526960224183 lpclm = -3.01910401042172e-05 wpclm = -3.68321342998292e-06 ppclm = 2.8902124220088e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.36784249985561e-05 lalpha0 = -1.0093911587572e-10 walpha0 = -1.23142596585178e-11 palpha0 = 9.66298231407536e-17   alpha1 = 0.0   beta0 = 18.7304132421031 lbeta0 = 6.46245339910028e-05 wbeta0 = 7.8839930880288e-06 pbeta0 = -6.18655833858588e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.402088621315792 lkt1 = 7.34369704443231e-08 wkt1 = 8.95908305457852e-09 pkt1 = -7.03017993021124e-14   kt2 = -0.019151   at = 571137.95921064 lat = -3.30466366999446 wat = -0.403158737456019 pat = 3.16358096859506e-6   ute = -1.33715518368426 lute = 1.32186546799778e-06 wute = 1.61263494982408e-07 pute = -1.26543238743803e-12   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.66 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.827662107734035+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.8060707516346e-07 wvth0 = -2.355816275876e-08 pvth0 = 1.84860573353712e-13   k1 = 0.88325   k2 = -0.0430122068799479 lk2 = 4.75308175860547e-08 wk2 = 3.97003492488122e-09 pk2 = -3.1152808475054e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 82241.0566868009 lvsat = 0.232733312953468 wvsat = 0.0283927437052721 pvsat = -2.22797462356858e-7   ua = -1.45894919862197e-10 lua = -2.03117674026134e-17 wua = -3.46964537756165e-18 pua = 2.72262587026913e-23   ub = 1.86433767298517e-18 lub = -6.39197219507186e-25 wub = -1.15811136251045e-25 pub = 9.08768364806048e-31   uc = 6.4498693309385e-11 luc = -9.30079184610372e-17 wuc = -1.13466781266206e-17 puc = 8.90372244060986e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0385865265269101 lu0 = -2.54136623252653e-10 wu0 = -2.4545136207377e-10 pu0 = 1.92605340187379e-15   a0 = 0.278738224445371 la0 = 6.61520455306864e-06 wa0 = 8.09729531924008e-07 pa0 = -6.35393630079425e-12   keta = -0.0175279297056782 lketa = -3.38210612585589e-08 wketa = -4.12606477331661e-09 pketa = 3.23771725113085e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.122727218075309 lags = 2.84347166352306e-07 wags = 2.47553467043509e-08 pags = -1.94254859014187e-13   b0 = -8.24430104923184e-08 lb0 = 9.05353939069076e-13 wb0 = 1.1045037785238e-13 pb0 = -8.66702568702339e-19   b1 = 9.31018719637085e-10 lb1 = -7.30569085873013e-15 wb1 = -8.91271668458339e-16 pb1 = 6.99379630458923e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.29282921115257+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.64017082364525e-06 wnfactor = -1.37848073108532e-07 pnfactor = 1.08169189980963e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.20949109728548 lpclm = 1.75559919183238e-05 wpclm = 2.14177666576017e-06 ppclm = -1.68064915113467e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.68995478935241e-05 lalpha0 = -2.04685082136813e-10 walpha0 = -1.65797994205557e-11 palpha0 = 1.30101453935908e-16   alpha1 = 0.0   beta0 = 27.6155554612656 lbeta0 = -5.09705261077438e-06 wbeta0 = -1.65667752261952e-06 pbeta0 = 1.29999253265102e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.394653493 lkt1 = 1.50936226420967e-8   kt2 = -0.019151   at = 310212.19447376 lat = -1.25718284706487 wat = -0.0520967774408662 pat = 4.08802683223593e-7   ute = -1.07074385694723 lute = -7.68660483149066e-07 wute = -9.37741993935594e-08 pute = 7.35844829802469e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.67 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.783127543335898+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.28322940773043e-09 wvth0 = 2.33971489419115e-08 pvth0 = 4.22414661559106e-15   k1 = 0.88325   k2 = -0.0335159618089194 lk2 = 1.09988957452391e-08 wk2 = -4.67071039579452e-09 pk2 = 2.08801780315119e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 175585.299273774 lvsat = -0.126360681459223 wvsat = -0.0592867187271747 pvsat = 1.14504202108291e-7   ua = -1.50332461453423e-10 lua = -3.24060702675122e-18 wua = 2.52761895885033e-18 pua = 4.15486676221488e-24   ub = 1.7341011811515e-18 lub = -1.38179258733952e-25 wub = 1.47580900263301e-25 pub = -1.04497112176135e-31   uc = -6.21897020841541e-12 luc = 1.79041943044652e-16 wuc = 4.47166979961739e-17 puc = -1.26637798651026e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0376550051046129 lu0 = 3.32941324702509e-09 wu0 = -2.06215456110547e-10 pu0 = 1.77511342093609e-15   a0 = 1.64687370831383 la0 = 1.35200650052344e-06 wa0 = -5.05397128771628e-07 pa0 = -1.29466244887138e-12   keta = -0.026319503488 wketa = 4.29017914109029e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.223964471257101 lags = -1.05111129316503e-07 wags = -4.50657552359174e-08 pags = 7.43459426545973e-14   b0 = 2.43480424583578e-07 lb0 = -3.48468952739807e-13 wb0 = -2.01558733933256e-13 pb0 = 3.3359211620944e-19   b1 = 3.95488682281792e-12 lb1 = -3.73928927278731e-15 wb1 = -3.78604479457858e-18 pb1 = 3.57965153515347e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.85938566910202+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.72804144136232e-08 wnfactor = 1.71469837253066e-07 pnfactor = -1.08249770900697e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.35407942736 wpclm = -2.22696590604715e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.72268081647873e-05 lalpha0 = -9.05344678187187e-11 walpha0 = 5.93567098580651e-13 palpha0 = 6.40357533639223e-17   alpha1 = 0.0   beta0 = 27.5907172603235 lbeta0 = -5.00150039948517e-06 wbeta0 = -8.28684015101206e-07 pbeta0 = 9.8146458949964e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352873999999 lkt1 = 6.39479635577644e-8   kt2 = -0.019151   at = -50370.2989475199 lat = 0.129972956971884 wat = 0.104193554881732 pat = -1.92444037156791e-7   ute = -1.36461228610554 lute = 3.61847249664919e-07 wute = 1.87548398787119e-07 pute = -3.46399266882225e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.68 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.748498513430697+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.46761040207576e-08 wvth0 = 4.75828761721818e-08 pvth0 = -4.04465529785376e-14   k1 = 0.88325   k2 = -0.0310810156928808 lk2 = 6.50158435816149e-09 wk2 = -7.24298188311797e-09 pk2 = 6.83896722843677e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 104171.262621021 lvsat = 0.00554004444189937 wvsat = 0.00752588045964708 pvsat = -8.89773321338037e-9   ua = -1.42038588355899e-10 lua = -1.85592745236559e-17 wua = -3.23207861155341e-18 pua = 1.47929475389847e-23   ub = 1.75208311881612e-18 lub = -1.71391645853385e-25 wub = 4.03519221383422e-26 pub = 9.35533092149692e-32   uc = 1.53846093695453e-10 luc = -1.16595989074899e-16 wuc = -6.84986022235435e-17 puc = 8.24692758405883e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0390291042895199 lu0 = 7.91471289890553e-10 wu0 = 1.72209339651345e-10 pu0 = 1.07616812111094e-15   a0 = 3.46649745652067 la0 = -2.00881308768212e-06 wa0 = -2.24455177900579e-06 pa0 = 1.91753184194601e-12   keta = -0.0395828837092872 lketa = 2.44972775813943e-08 wketa = 7.92390081108583e-09 pketa = -6.71143305237834e-15   a1 = 0.0   a2 = 0.65972622   ags = 0.164988942332243 lags = 3.8158469503038e-09 wags = -3.35189182313404e-09 pags = -2.69897907472542e-15   b0 = -1.16418536551211e-09 lb0 = 1.03386216811623e-13 wb0 = 3.26415083278876e-14 pb0 = -9.89724524435009e-20   b1 = -3.3665937946422e-09 lb1 = 2.48606695419703e-15 wb1 = 3.22286717236133e-15 pb1 = -2.37993178378845e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.846788179556614+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.054780123913e-08 wnfactor = 1.47225325395055e-07 pnfactor = -6.34704969221129e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 5.9402597473732 lpclm = -4.7766388445399e-06 wpclm = -4.70273701583834e-06 ppclm = 4.5727145789888e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -6.68336329063158e-05 lalpha0 = 8.31938499934336e-11 walpha0 = 6.71232695517004e-11 palpha0 = -5.88436756511555e-17   alpha1 = 0.0   beta0 = 15.9054108582907 lbeta0 = 1.65810969307798e-05 wbeta0 = 8.28407812068064e-06 pbeta0 = -7.01649819112279e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16612.056 lat = 0.00625748513678401   ute = -1.73263548352947 lute = 1.04158094298215e-06 wute = 4.76696567566331e-07 pute = -8.80451886543067e-13   ua1 = 3.0044e-9   ub1 = -4.49406467598122e-18 lub1 = 1.36965957463186e-24 wub1 = 3.44790635732529e-25 pub1 = -6.36823477129079e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.69 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.760572682771906+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.44494516271253e-08 wvth0 = 3.51913251270082e-08 pvth0 = -2.99510827249885e-14   k1 = 0.88325   k2 = -0.0381123220051035 lk2 = 1.24570023663257e-08 wk2 = 4.51996598779804e-09 pk2 = -3.12408493695884e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 145884.657563996 lvsat = -0.029790617087271 wvsat = -0.0365381039211359 pvsat = 2.84238446613614e-8   ua = -2.24590293099842e-10 lua = 5.13608636705981e-17 wua = 5.68486834009032e-17 pua = -3.60946167548978e-23   ub = 1.20227278027029e-18 lub = 2.94290013550194e-25 wub = 1.77616898961558e-25 pub = -2.2708204444615e-32   uc = -1.97096944797034e-10 luc = 1.80647851325699e-16 wuc = 1.72770417166443e-16 puc = -1.21882205816459e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0400720309300254 lu0 = -9.1872973644637e-11 wu0 = 9.45063890352703e-10 pu0 = 4.21571136630647e-16   a0 = 1.00607018913251 la0 = 7.51343618139148e-08 wa0 = 8.21395442650628e-08 pa0 = -5.31431351858763e-14   keta = 0.0459272576167633 lketa = -4.79286149797919e-08 wketa = -5.41714344145884e-08 pketa = 4.58824465490746e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.199398323802604 lags = -2.53284174237516e-08 wags = -2.76899226121721e-08 pags = 1.79149922711589e-14   b0 = 4.05464890838146e-07 lb0 = -2.41022917925809e-13 wb0 = -3.56627759354484e-13 pb0 = 2.3073316751372e-19   b1 = -1.82695428775892e-09 lb1 = 1.18201384681999e-15 wb1 = 1.74895795530592e-15 pb1 = -1.13155131167156e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.918095599563536+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.84858520285322e-09 wnfactor = 2.83926457949319e-08 pnfactor = 3.71791190416726e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.34582353252942 lpclm = 1.3945716883717e-06 wpclm = 2.27228879667868e-06 ppclm = -1.33503463385174e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.699649258132e-05 lalpha0 = 3.72104732716281e-12 walpha0 = -8.92215745020952e-12 palpha0 = 5.5657363834842e-18   alpha1 = 0.0   beta0 = 30.7007734599999 lbeta0 = 4.04963194220842e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37919986 lkt1 = 5.47988084196013e-9   kt2 = -0.019151   at = 7825.35000000003 lat = 0.0136997021049   ute = 1.90459592964732 lute = -2.0391031427388e-06 wute = -2.38348283783165e-06 pute = 1.54208002731735e-12   ua1 = 6.21571501100001e-09 lua1 = -2.71993885590685e-15   ub1 = -6.35699552909388e-18 lub1 = 2.94753592618633e-24 wub1 = -1.72395317866264e-24 pub1 = 1.11537357125023e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.70 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784585564548125+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.89134532982541e-08 wvth0 = 4.03710171731757e-09 pvth0 = -9.79473633804753e-15   k1 = 0.88325   k2 = -0.00486654972190897 lk2 = -9.05254686008918e-09 wk2 = -1.22868180146204e-08 pk2 = 7.74966901762981e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 158428.664364397 lvsat = -0.0379064138710359 wvsat = -0.0403117862015888 pvsat = 3.08653642652625e-8   ua = -1.381368010052e-10 lua = -4.57333536574588e-18 wua = -5.65317059802917e-18 pua = 4.34320775645533e-24   ub = 3.5381646889732e-19 lub = 8.4322936862015e-25 wub = 6.09037663591721e-25 pub = -3.01831399269625e-31   uc = 1.68012270954224e-10 luc = -5.55726997363444e-17 wuc = -8.39607413282077e-17 puc = 4.42192594933613e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0312457234593309 lu0 = 5.61862439159009e-09 wu0 = 4.33856890067818e-09 pu0 = -1.77397909597983e-15   a0 = 1.1222   keta = -0.0281525756096 wketa = 1.6745782571675e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.986644924627466+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.41990388286629e-08 wnfactor = -5.84804908747577e-09 pnfactor = 5.93323692608651e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -5.34786189557032 lpclm = 3.98383448072208e-06 wpclm = 4.56409011083205e-06 ppclm = -2.81779799889057e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 6.00867813961969e-05 lalpha0 = -1.76879062720192e-11 walpha0 = 7.63924004726584e-13 palpha0 = -7.01022712719134e-19   alpha1 = 0.0   beta0 = 34.6836712294464 lbeta0 = 1.47275284594539e-06 wbeta0 = 2.17914774268109e-06 pbeta0 = -1.40987808144629e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.71 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.918523003111869+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.09547066155973e-08 wvth0 = -3.58069967100407e-08 pvth0 = 8.01501784160418e-15   k1 = 0.88325   k2 = -0.00466861939409946 lk2 = -9.14101894559545e-09 wk2 = -2.62252364969873e-09 pk2 = 3.42986473663092e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -42309.1992762547 lvsat = 0.0518206008462448 wvsat = 0.105894593690872 pvsat = -3.44868406573491e-8   ua = -1.60323066114063e-10 lua = 5.34361453020438e-18 wua = 1.66160636967771e-19 pua = 1.742048165049e-24   ub = 2.3376039370374e-18 lub = -4.34958566139143e-26 wub = -1.08025815360265e-24 pub = 4.53260180874815e-31   uc = -4.74331287962072e-11 luc = 4.0728377716502e-17 wuc = 1.45297367099394e-16 puc = -5.82559053602589e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0350017808810013 lu0 = 3.93971930890731e-09 wu0 = 4.47087993403154e-09 pu0 = -1.83312027553427e-15   a0 = 1.1222   keta = -0.0888493640143266 lketa = 2.71306146618751e-08 wketa = 7.4851303685827e-08 pketa = -2.59723544607304e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.423001150890602+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.97741837018881e-07 wnfactor = 3.83078284766574e-07 pnfactor = -1.14512257003221e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 11.4760747066868 lpclm = -3.53622964537445e-06 wpclm = -7.77713616610197e-06 ppclm = 2.69855736973106e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.15019733514135e-05 lalpha0 = -9.38075726331355e-12 walpha0 = -3.59559377542387e-12 palpha0 = 1.24762070175923e-18   alpha1 = 0.0   beta0 = 41.5126575411072 lbeta0 = -1.57970842955862e-06 wbeta0 = -4.35829548536229e-06 pbeta0 = 1.51226751728388e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4401272 lkt1 = 3.10195768392001e-8   kt2 = -0.019151   at = 29739.22944 lat = 0.00387124318953216   ute = -1.841439118 lute = 2.42417992998348e-7   ua1 = -1.432830022e-09 lua1 = 1.53965669641369e-15   ub1 = -4.30134779151005e-18 lub1 = 1.11753106073591e-24 wub1 = 2.25456338799332e-24 pub1 = -1.00775827054558e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.72 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.815346+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.036493   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 101000.0   ua = -1.460743e-10   ub = 1.86843e-18   uc = 5.7002e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03888129   a0 = 0.80798   keta = -0.020254   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -9.469e-9   b1 = 3.4216e-10   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.06912+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.20557   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8066e-5   alpha1 = 0.0   beta0 = 28.726   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.39073   kt2 = -0.019151   at = 60000.0   ute = -1.1327   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.73 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.822342895849999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.38867293978393e-7   k1 = 0.88325   k2 = -0.036190891039 lk2 = -5.9959523194417e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93872.3210499999 lvsat = 0.141462944333146   ua = -1.4449895216895e-10 lua = -3.12659063479796e-17   ub = 1.924372471025e-18 lub = -1.11028943923858e-24   uc = 5.98504559179999e-11 luc = -5.65332647261631e-17 wuc = 9.86076131526265e-32   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.039095218455825 lu0 = -4.24583506776034e-9   a0 = 0.602792354193635 la0 = 4.07235633369179e-6   keta = -0.019218197848 lketa = -2.05575508095147e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16109113150765 lags = -1.66939252564876e-8   b0 = -3.7196325031e-08 lb0 = 5.50303831707707e-13 pb0 = -3.85185988877447e-34   b1 = 5.65903727479999e-10 lb1 = -4.44063862688337e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.059513981305+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.90650518555374e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.332098941565 lpclm = 1.06711079558754e-05 ppclm = 6.46234853557053e-27   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.62683862904999e-05 lalpha0 = 3.56772141258551e-11   alpha1 = 0.0   beta0 = 29.87689128 lbeta0 = -2.28417231216815e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.389422169000001 lkt1 = -2.59565035473609e-8   kt2 = -0.019151   at = 1147.60499999998 lat = 1.16804265963147 pat = -8.470329472543e-22   ute = -1.109159042 lute = -4.67217063852604e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.74 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.794355312449998+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.07508811352095e-8   k1 = 0.88325   k2 = -0.0373993268830001 lk2 = 3.48662683032398e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 122383.03685 lvsat = -0.0822602433994337   ua = -1.50800343493151e-10 lua = 1.81810231535397e-17   ub = 1.70060258692499e-18 lub = 6.45629708515729e-25   uc = 4.84566322459998e-11 luc = 3.28739101144899e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.038239504632525 lu0 = 2.46893932368227e-9   a0 = 1.42354293741908 la0 = -2.36806200237006e-6   keta = -0.0233614064559999 lketa = 1.19541491325417e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.15772660547705 lags = 9.70746340226924e-9   b0 = 7.37129750930001e-08 lb0 = -3.1999989363512e-13   b1 = -3.29071182440001e-10 lb1 = 2.58221696161013e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.097938056085+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.10862658306209e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.818576824695 lpclm = -6.20521467250612e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.34588411285001e-05 lalpha0 = -2.07461843215636e-11   alpha1 = 0.0   beta0 = 25.2733261600001 lbeta0 = 1.32823879250466e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.394653493 lkt1 = 1.50936226421018e-8   kt2 = -0.019151   at = 236557.185 lat = -0.67921301889441   ute = -1.203322874 lute = 2.71685207557778e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.75 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.816206695475998+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.3110834464373e-9   k1 = 0.88325   k2 = -0.0401194646617 lk2 = 1.39509587830546e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 91765.0699999998 lvsat = 0.0355266464209798   ua = -1.467588853609e-10 lua = 2.63359029918728e-18   ub = 1.94275271663999e-18 lub = -2.85918450396042e-25   uc = 5.7002e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0373634553750601 lu0 = 5.83908855245938e-9   a0 = 0.932337567379999 la0 = -4.78401820704915e-7   keta = -0.020254   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -4.14855788170001e-08 lb0 = 1.23167330476895e-13   b1 = -1.39786586000016e-12 lb1 = 1.3216623001533e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.1018116522+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.25764328330265e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.20557   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8066e-5   alpha1 = 0.0   beta0 = 26.419114486 lbeta0 = 8.8745562759607e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874000001 lkt1 = 6.39479635577652e-8   kt2 = -0.019151   at = 96939.72 lat = -0.142106585683921   ute = -1.099454252 lute = -1.2789592711553e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.76 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.815771718557997+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.50768716856465e-9   k1 = 0.88325   k2 = -0.0413212248848001 lk2 = 1.61705930904771e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 114811.437 lvsat = -0.00703967077888157   ua = -1.46608137423e-10 lua = 2.35516096835672e-18   ub = 1.80913311986001e-18 lub = -3.91249258177438e-26   uc = 5.7002e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0392725757894201 lu0 = 2.3129698748224e-9   a0 = 0.293124924320004 la0 = 7.02214982049902e-7   keta = -0.028379983684 lketa = 1.50085781005764e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 4.4984745974e-08 lb0 = -3.65421488275344e-14   b1 = 1.1899320362e-09 lb1 = -8.78707350332889e-16 wb1 = 1.57772181044202e-30   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.0549369993+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.9187500669109e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.70852270078 lpclm = 1.68831642104285e-06 wpclm = -4.2351647362715e-22 ppclm = -8.07793566946316e-28   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8066e-5   alpha1 = 0.0   beta0 = 27.6175336120001 lbeta0 = 6.66109292810665e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16612.056 lat = 0.00625748513678404   ute = -1.0586765186 lute = -2.03211829817062e-7   ua1 = 3.0044e-9   ub1 = -4.0065958e-18 lub1 = 4.69311385258809e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.77 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.810326573760008+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.10427424330385e-9   k1 = 0.88325   k2 = -0.0317219432906002 lk2 = 8.04013597013201e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 94226.6755800014 lvsat = 0.0103953339571978   ua = -1.44216985572001e-10 lua = 3.29888826685926e-19   ub = 1.45338954830003e-18 lub = 2.62184898883581e-25   uc = 4.71678128000005e-11 luc = 8.32941887977963e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0414081728800006 lu0 = 5.04149037460191e-10   a0 = 1.1222   keta = -0.030660925204 lketa = 1.69405036348352e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -9.87394435599997e-08 lb0 = 8.51902275691101e-14 wb0 = -2.52435489670724e-29 pb0 = -2.40741243048404e-35   b1 = 6.457421264e-10 lb1 = -4.17786115391031e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.9582374413+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.27156711630829e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.86676390700001 lpclm = -4.92915281734296e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.43822461000003e-05 lalpha0 = 1.15899479807454e-11   alpha1 = 0.0   beta0 = 30.7007734600006 lbeta0 = 4.04963194220831e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37919986 lkt1 = 5.47988084195843e-9   kt2 = -0.019151   at = 7825.35000000033 lat = 0.0136997021049   ute = -1.465198895 lute = 1.41106931680474e-7   ua1 = 6.21571501100003e-09 lua1 = -2.71993885590685e-15   ub1 = -8.79433990900001e-18 lub1 = 4.52446361716427e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.78 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.790293264329996+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.50655449781897e-8   k1 = 0.88325   k2 = -0.0222377911253999 lk2 = 1.90402229737804e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 101435.407959001 lvsat = 0.00573138503023829   ua = -1.46129317133999e-10 lua = 1.56714057465822e-18   ub = 1.21488076280001e-18 lub = 4.16496743979082e-25   uc = 4.93076312099999e-11 luc = 6.94498632596707e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0373796409332998 lu0 = 3.11055280752794e-9   a0 = 1.1222   keta = -0.0044772   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.978376887099991+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.96857316827161e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.1049   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 6.11668257400001e-05 lalpha0 = -1.86790200622196e-11   alpha1 = 0.0   beta0 = 37.7645748 lbeta0 = -5.20548631552788e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.65799999982 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909577e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.79 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.867898668719995+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.96229843084794e-8   k1 = 0.88325   k2 = -0.00837637280519976 lk2 = -4.29183763189488e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 107405.767457999 lvsat = 0.00306271791921864   ua = -1.60088146337999e-10 lua = 7.80654180523744e-18   ub = 8.10322818199962e-19 lub = 5.97328481404056e-25   uc = 1.5798992184e-10 luc = -4.16344760335743e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0413227611809996 lu0 = 1.34803326048948e-9   a0 = 1.1222   keta = 0.016976250408 lketa = -9.58939198407031e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.964601535399993+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.58431210376995e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.480672185999993 lpclm = 2.79021093668606e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.641848246e-05 lalpha0 = -7.61685709286556e-12   alpha1 = 0.0   beta0 = 35.3508503999997 lbeta0 = 5.58352383105555e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.440127199999999 lkt1 = 3.10195768392005e-8   kt2 = -0.019151   at = 29739.2294399999 lat = 0.00387124318953214   ute = -1.841439118 lute = 2.42417992998347e-7   ua1 = -1.43283002200002e-09 lua1 = 1.53965669641369e-15   ub1 = -1.11382073399998e-18 lub1 = -3.07248908592274e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.80 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.832257483571428+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.11160534433686e-8   k1 = 0.88325   k2 = -0.0330442701271429 wk2 = -2.26687773526798e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 63673.4585714286 wvsat = 0.0245350342933314   ua = -3.52541684444286e-10 wua = 1.35712663534305e-16   ub = 1.81650702908571e-18 wub = 3.41293841657275e-26   uc = 2.85462391571429e-11 wuc = 1.87041992480967e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0352246229932857 wu0 = 2.40355647684935e-9   a0 = 0.409084592285715 wa0 = 2.62197142653862e-7   keta = -0.0274821432571429 wketa = 4.75111638806606e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -6.46794016171429e-08 wb0 = 3.62902386661609e-14   b1 = 1.68862402385714e-09 wb1 = -8.85041574593491e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.797916399714286+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.78264296096602e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.191142411428571 wpclm = 2.60762241731291e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.54585226857143e-05 walpha0 = 8.28699569849852e-12   alpha1 = 0.0   beta0 = 34.7332823714286 wbeta0 = -3.94863476099897e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.394772585714286 wkt1 = 2.65722393068575e-9   kt2 = -0.019151   at = -209505.714285714 wat = 0.177148262045714   ute = -1.25909818 wute = 8.308253489944e-8   ua1 = 3.0044e-9   ub1 = -4.15702807714286e-18 wub1 = 2.65899541330616e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.81 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.851973184596813+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.91297242230995e-07 wvth0 = -1.94762258355904e-08 pvth0 = 1.65924224426014e-13   k1 = 0.88325   k2 = -0.0327055045016496 lk2 = -6.72347662644641e-09 wk2 = -2.29097245409273e-09 pk2 = 4.78207547188775e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 46941.0285883336 lvsat = 0.332088303620467 wvsat = 0.030848313985393 pvsat = -1.25299573662431e-7   ua = -3.47629082155654e-10 lua = -9.75003488460429e-17 wua = 1.335190594813e-16 pua = 4.35364289295166e-23   ub = 1.95948264318767e-18 lub = -2.83763501142286e-24 wub = -2.30781970438986e-26 pub = 1.13539806336131e-30   uc = 3.52330708091027e-11 luc = -1.32713454180803e-16 wuc = 1.61812041711591e-17 puc = 5.00738479700505e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0356938704043253 lu0 = -9.31314679743948e-09 wu0 = 2.23573328503515e-09 pu0 = 3.33078453841184e-15   a0 = -0.248004933028505 la0 = 1.30412466096579e-05 wa0 = 5.59235863269414e-07 pa0 = -5.89532332951477e-12   keta = -0.0250505681109757 lketa = -4.82594378839284e-08 wketa = 3.833663632816e-09 pketa = 1.82086719891092e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.162224580246537 lags = -3.91894665088992e-08 wags = -7.45024923660423e-10 pags = 1.478649922954e-14   b0 = -1.27051504209426e-07 lb0 = 1.23789824693961e-12 wb0 = 5.9062528115413e-14 pb0 = -4.51961309887254e-19   b1 = 3.09867786769911e-09 lb1 = -2.79853188979778e-14 wb1 = -1.66481270455914e-15 pb1 = 1.54761066996325e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.678137718480949+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.37724580953649e-06 wnfactor = 2.50681668564351e-07 pnfactor = -1.4372665775242e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.45333561372217 lpclm = 2.50507308152162e-05 wpclm = 7.36997834502284e-07 ppclm = -9.45184114242759e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -3.41704329648427e-06 lalpha0 = 3.74623093790771e-10 walpha0 = 1.95124703509615e-11 palpha0 = -2.22791838270787e-16   alpha1 = 0.0   beta0 = 38.3258952214016 lbeta0 = -7.13025369368351e-05 wbeta0 = -5.55359788271481e-06 pbeta0 = 3.18536806072107e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.404919962368436 lkt1 = 2.01394842391642e-07 wkt1 = 1.01868235634197e-08 pkt1 = -1.49439858496477e-13   kt2 = -0.019151   at = -407582.940774614 lat = 3.93123594104403 wat = 0.26866185758202 pat = -1.81626904941873e-6   ute = -1.27247823743915 lute = 2.65553812673907e-07 wute = 1.07351013715714e-07 pute = -4.81656159307878e-13   ua1 = 3.0044e-9   ub1 = -4.42155525697177e-18 lub1 = 5.25006723468385e-24 wub1 = 4.39775372849598e-25 pub1 = -3.45091119389558e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.82 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.779993334987307+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.73527629936902e-07 wvth0 = 9.44024268204759e-09 pvth0 = -6.09828992013334e-14   k1 = 0.88325   k2 = -0.0309894810951741 lk2 = -2.01890882727317e-08 wk2 = -4.21324291510426e-09 pk2 = 1.55622369429599e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 106094.863197385 lvsat = -0.132091008403075 wvsat = 0.0107063468472531 pvsat = 3.27541604830133e-8   ua = -3.64924305243833e-10 lua = 3.8215024593779e-17 wua = 1.40745393050418e-16 pua = -1.31685094186813e-23   ub = 1.37602910913205e-18 lub = 1.74071670196208e-24 wub = 2.13344743541129e-25 pub = -7.1980944148823e-31   uc = -2.34122333759176e-11 luc = 3.27475426724792e-16 wuc = 4.72399803242114e-17 puc = -1.93643933680085e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.034091110315903 lu0 = 3.2636891777697e-09 wu0 = 2.72677277147021e-09 pu0 = -5.22395437091304e-16   a0 = 2.12237521281808 la0 = -5.55909320947811e-06 wa0 = -4.59348045277962e-07 pa0 = 2.09749034068177e-12   keta = -0.0422805980326565 lketa = 8.69443656910825e-08 wketa = 1.24357359768689e-08 pketa = -4.92916692656614e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.154326259260389 lags = 2.2788547692915e-08 wags = 2.23507477098132e-09 pags = -8.59830135291833e-15   b0 = 1.0295623985535e-07 lb0 = -5.66969300628268e-13 wb0 = -1.92218318744106e-14 pb0 = 1.62334966971852e-19   b1 = -1.72586787294579e-09 lb1 = 9.87282398522246e-15 wb1 = 9.18125639042982e-16 pb1 = -4.79217432147657e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.918766040547808+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.89038735074364e-07 wnfactor = 1.17771199188721e-07 pnfactor = -3.94319985080197e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.59543719545222 lpclm = -1.45669187355559e-05 wpclm = -1.16794453658169e-06 ppclm = 5.49621497427513e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.25614800405186e-05 lalpha0 = 1.38302648646363e-11 walpha0 = -5.9832373779811e-12 palpha0 = -2.27273766616827e-17   alpha1 = 0.0   beta0 = 26.6303483727345 lbeta0 = 2.04722554470001e-05 wbeta0 = -8.91981556608063e-07 pbeta0 = -4.72595744112048e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.3682183984135 lkt1 = -8.66018161408421e-08 wkt1 = -1.73759991524631e-08 pkt1 = 6.68452254755371e-14   kt2 = -0.019151   at = 151449.405481129 lat = -0.455483053571939 wat = 0.0559420243399903 pat = -1.47059496046183e-7   ute = -1.34052101490394 lute = 7.99484534841229e-07 wute = 9.01814356012838e-08 pute = -3.46926720218041e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.83 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.817508020056495+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.92091616813264e-08 wvth0 = -8.55371057356266e-10 pvth0 = -2.1375817284439e-14   k1 = 0.88325   k2 = -0.0386788995053266 lk2 = 9.39199669926725e-09 wk2 = -9.46895001805469e-10 pk2 = 2.99664224937016e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 47590.5015638286 lvsat = 0.0929744517401534 wvsat = 0.029036297229643 pvsat = -3.77609020187352e-8   ua = -4.4989353570134e-10 lua = 3.65090464594581e-16 wua = 1.99252830745974e-16 pua = -2.38245803129357e-22   ub = 1.96540041386479e-18 lub = -5.26586456146503e-25 wub = -1.48865125674326e-26 pub = 1.58193005523819e-31   uc = 7.07923445349065e-11 luc = -3.49282656340574e-17 wuc = -9.06450378555032e-18 puc = 2.2958628427391e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.033705531424903 lu0 = 4.7470057733419e-09 wu0 = 2.40438267582977e-09 pu0 = 7.17834747376131e-16   a0 = 0.848596328847925 la0 = -6.58883675749321e-07 wa0 = 5.50437860170416e-08 pa0 = 1.18632167175526e-13   keta = -0.0196799528285714 wketa = -3.77325798157371e-10   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -1.13154982748388e-07 lb0 = 2.64407547171193e-13 wb0 = 4.71088725593325e-14 pb0 = -9.28383243548954e-20   b1 = 2.98189469930341e-09 lb1 = -8.23787272154421e-15 wb1 = -1.96094206942243e-15 pb1 = 6.28355884604194e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.04780542651803+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.37397620167237e-09 wnfactor = 3.54987241905654e-08 pnfactor = -7.78189255769431e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.191142411428572 wpclm = 2.60762241731291e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.77407345388657e-05 lalpha0 = -6.09425468094231e-12 walpha0 = -1.29323604102728e-11 palpha0 = 4.00580235582084e-18   alpha1 = 0.0   beta0 = 31.0052633768946 lbeta0 = 3.6420186748061e-06 wbeta0 = -3.01451235517615e-06 pbeta0 = 3.43938882553978e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407352874 lkt1 = 6.3947963557764e-8   kt2 = -0.019151   at = 45100.4845111428 lat = -0.0463602434852978 wat = 0.0340743442007097 pat = -6.2934836697892e-8   ute = -1.099454252 lute = -1.27895927115529e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.84 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.829085401407077+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.82590041014192e-09 wvth0 = -8.75119024616069e-09 pvth0 = -6.79234978418559e-15   k1 = 0.88325   k2 = -0.0417413366630875 lk2 = 1.50482752555314e-08 wk2 = 2.76142832762627e-10 pk2 = 7.3770849145257e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110357.510508373 lvsat = -0.0229553350422947 wvsat = 0.00292760151435845 pvsat = 1.04614934456553e-8   ua = -2.52104809188851e-10 lua = -2.22544231815205e-19 wua = 6.93438063250681e-17 pua = 1.69434624971485e-24   ub = 1.62893314065499e-18 lub = 9.48638869301743e-26 wub = 1.18446887931287e-25 pub = -8.8071918529708e-32   uc = 5.18813914285715e-11 wuc = 3.36581697886857e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0353558109903611 lu0 = 1.69896251985489e-09 wu0 = 2.57452083653984e-09 pu0 = 4.03591946478937e-16   a0 = -0.0420258259158071 la0 = 9.86082975389126e-07 wa0 = 2.20297269335998e-07 pa0 = -1.8658870296582e-13   keta = -0.0273197265950318 lketa = 1.41105551898196e-08 wketa = -6.96915466635492e-10 pketa = 5.9027764342373e-16   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 1.34440158804117e-07 lb0 = -1.928972129443e-13 wb0 = -5.87997584965383e-14 pb0 = 1.02773434484463e-19   b1 = -2.38066650860852e-09 lb1 = 1.66670275361221e-15 wb1 = 2.346982988291e-15 pb1 = -1.67311842460395e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05322855509024+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.73904187507408e-08 wnfactor = 1.12297404663148e-09 pnfactor = -1.43273963215992e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.61073363915291 lpclm = 2.62196512332967e-06 wpclm = 5.93030467480022e-07 ppclm = -6.13694761202744e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.27896513533338e-05 lalpha0 = 3.05032664757061e-12 walpha0 = -9.67797382375713e-12 palpha0 = -2.00500410806135e-18   alpha1 = 0.0   beta0 = 27.480612829331 lbeta0 = 1.01519988910485e-05 wbeta0 = 8.99991258146129e-08 pbeta0 = -2.29460041668942e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16612.056 lat = 0.00625748513678399   ute = -1.0586765186 lute = -2.0321182981706e-7   ua1 = 3.0044e-9   ub1 = -4.34899715038e-18 lub1 = 1.10172188579175e-24 wub1 = 2.25063146815577e-25 pub1 = -4.15688481284316e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.85 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.846873715214004+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.24055234793259e-09 wvth0 = -2.40227284548495e-08 pvth0 = 6.14242927703873e-15   k1 = 0.88325   k2 = -0.0329816042356541 lk2 = 7.62890452574929e-09 wk2 = 8.27985216471629e-10 pk2 = 2.70305718244409e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 29396.7233320462 lvsat = 0.0456173182450336 wvsat = 0.042613246252198 pvsat = -2.31516920482685e-8   ua = -3.96643780399752e-10 lua = 1.22199940838221e-16 wua = 1.6592215165464e-16 pua = -8.01061601475981e-23   ub = 1.18042753089611e-18 lub = 4.74741859317412e-25 wub = 1.79420117735719e-25 pub = -1.39715390548845e-31   uc = -8.30981904078168e-12 luc = 5.09811125905954e-17 wuc = 3.64658912300005e-17 puc = -2.80352994896692e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.036405537465047 lu0 = 8.09858891966543e-10 wu0 = 3.28827227933191e-09 pu0 = -2.00945533045761e-16   a0 = 1.1222   keta = -0.0576127433713958 lketa = 3.9768316297165e-08 wketa = 1.77156456959746e-08 pketa = -1.50049038854507e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -5.01677352687184e-07 lb0 = 3.4588541364367e-13 wb0 = 2.64854311172571e-13 pb0 = -1.71357031368297e-19   b1 = -1.74844224924042e-09 lb1 = 1.13121765706706e-15 wb1 = 1.57371654358345e-15 pb1 = -1.01817257166688e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.994077200958829+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.2709950079602e-08 wnfactor = -2.35577607418257e-08 pnfactor = 6.57684051393712e-15   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.85108489207984 lpclm = -1.15713270716504e-06 wpclm = -6.47002058060861e-07 ppclm = 4.36595427475026e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -5.9122602907048e-06 lalpha0 = 4.43001639833082e-11 walpha0 = 1.33397414066613e-11 palpha0 = -2.15006866602126e-17   alpha1 = 0.0   beta0 = 28.2425760765917 lbeta0 = 9.50662668810411e-06 wbeta0 = 1.61579280569333e-06 pbeta0 = -3.58692630243518e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37919986 lkt1 = 5.4798808419597e-9   kt2 = -0.019151   at = 7825.34999999998 lat = 0.0136997021049   ute = -1.465198895 lute = 1.41106931680469e-7   ua1 = 6.215715011e-09 lua1 = -2.71993885590685e-15   ub1 = -7.0823331571e-18 lub1 = 3.4168192167795e-24 wub1 = -1.12531573407788e-24 pub1 = 7.28063525528113e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.86 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.789731232828288+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.97298337608724e-08 wvth0 = 3.69427802327166e-10 pvth0 = -9.63895433116691e-15   k1 = 0.88325   k2 = -0.0158332461660316 lk2 = -3.46584306828355e-09 wk2 = -4.20975863815254e-09 pk2 = 3.52965546377229e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 70665.8444667377 lvsat = 0.0189167746385841 wvsat = 0.020225080239972 pvsat = -8.66686207268245e-9   ua = -2.08629357527063e-10 lua = 5.57241441511128e-19 wua = 4.10817765506832e-17 pua = 6.63814779410589e-25   ub = 1.04177962103697e-18 lub = 5.64445115925539e-25 wub = 1.13780765289976e-25 pub = -9.72476484673829e-32   uc = 4.52888040549381e-11 luc = 1.63035538283881e-17 wuc = 2.6416072396394e-18 puc = -6.15146128788146e-24   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0310799145172798 lu0 = 4.25546238045066e-09 wu0 = 4.14086057106141e-09 pu0 = -7.52558221558657e-16   a0 = 1.1222   keta = 0.00385429965142857 wketa = -5.47636137288122e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.876388909715295+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.08852626878092e-07 wnfactor = 6.70375134387851e-08 pnfactor = -5.20370335470799e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.36301031347283 lpclm = -8.41355287850399e-07 wpclm = -8.26965973928197e-07 ppclm = 5.5302956154637e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 0.000130334423973957 lalpha0 = -4.38495332823481e-11 walpha0 = -4.54644156599657e-11 palpha0 = 1.65447797036962e-17   alpha1 = 0.0   beta0 = 48.7431848163531 lbeta0 = -3.7569801579991e-06 wbeta0 = -7.21632819262896e-06 pbeta0 = 2.12733233378536e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 7991.658 lat = 0.013592103157212   ute = -1.13088364 lute = -7.51903578909594e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.87 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 7.6507e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 2.1346e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.894214847305843+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.69728791399921e-08 wvth0 = -1.72978347139033e-08 pvth0 = -1.74193532808731e-15   k1 = 0.88325   k2 = -0.000736395436463061 lk2 = -1.02139239884904e-08 wk2 = -5.02181824428971e-09 pk2 = 3.89263473888111e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 116726.587359479 lvsat = -0.00167173258407105 wvsat = -0.00612664948780173 pvsat = 3.11199219141619e-9   ua = -4.95477239471713e-10 lua = 1.28774228800423e-16 wua = 2.20453934029535e-16 pua = -7.95130284034315e-23   ub = 5.86438938249096e-19 lub = 7.67976026362156e-25 wub = 1.47160665362765e-25 pub = -1.12167996481319e-31   uc = 2.33612002116887e-10 luc = -6.78742791805303e-17 wuc = -4.97069983426402e-17 puc = 1.72476325269194e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0354333618312083 lu0 = 2.30953237938698e-09 wu0 = 3.87114930781284e-09 pu0 = -6.32001062844237e-16   a0 = 1.1222   keta = 0.0542168874399346 lketa = -2.25113716652331e-08 wketa = -2.44785686461868e-08 pketa = 8.49372062026579e-15   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.21328955460352+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.17372447779159e-08 wnfactor = -1.63464624526627e-07 pnfactor = 5.09941950935281e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.266942465191544 lpclm = 3.34196784873673e-07 wpclm = 4.91413091145411e-07 ppclm = -3.62674232346212e-14   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 9.38828309007499e-05 lalpha0 = -2.75561815009276e-11 walpha0 = -3.77717759448924e-11 palpha0 = 1.31062774480145e-17   alpha1 = 0.0   beta0 = 52.0593849032326 lbeta0 = -5.23927517003306e-06 wbeta0 = -1.09826533972508e-05 pbeta0 = 3.81082697169847e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.369991167667143 lkt1 = -3.30247709134448e-10 wkt1 = -4.61009751406457e-08 pkt1 = 2.06064904742167e-14   kt2 = -0.019151   at = 70436.8311350127 lat = -0.0143200150017147 wat = -0.0267508591749454 pat = 1.19572595391721e-8   ute = -2.56991870716394 lute = 5.68038170640383e-07 wute = 4.78835461794173e-07 pute = -2.14032747725531e-13   ua1 = -1.43283002200001e-09 lua1 = 1.5396566964137e-15   ub1 = -9.31132019306436e-18 lub1 = 3.35691858461706e-24 wub1 = 5.38828197443867e-24 pub1 = -2.40848660662645e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 2.75467857e-10   cgso = 2.75467857e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 4.49025e-11   cgdl = 4.49025e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 6.5995e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00084698656   mjs = 0.295   pbs = 0.72468   cjsws = 8.64309376e-11   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 5.47776e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__nfet_g5v0d10v5





















