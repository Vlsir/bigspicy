** Translated using xdm 2.6.0 on Nov_14_2022_16_05_13_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX_SLOPE=0.80e-2
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__tox2_slope=0.86e-2  ; for L>=4 and W<=0.75; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__tox3_slope=0.55e-2  ; for L>=4 and W>=3.0; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__tox4_slope=2.55e-2  ; for L<=0.6 and W<=3.0; HSpice Parser Retained (as a comment). Continuing.
.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__TOX_OFFSET=0.000
.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__NFACTOR_SLOPE=0.000
.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__VOFF_SLOPE=0.00375
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__voff2_slope=0.00850 ; for L>=4 and W=0.42; HSpice Parser Retained (as a comment). Continuing.
.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__LINT_SLOPE=3.0e-09
.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__LINT1_SLOPE=0.0e-09
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__wint_slope=0.0e-11  ; Not used; HSpice Parser Retained (as a comment). Continuing.
.PARAM SKY130_FD_PR__RF_NFET_G5V0D10V5__B_TOXE_SLOPE=.80e-2
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1= 2.05e-2 ; All W with L=0.5um; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope2= 1.00e-2 ; W=3 L=1 um All W with L=0.8um & L=0.6um; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope3= 0.67e-2 ; All W with L=4.0um; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_vth0_slope=0.000  ; All devices; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope=0.13  ; All devices; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope=0.12  ; All devices; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_lint_slope=0.0  ; All devices; HSpice Parser Retained (as a comment). Continuing.
* .param sky130_fd_pr__rf_nfet_g5v0d10v5__b_wint_slope=0.0  ; All devices; HSpice Parser Retained (as a comment). Continuing.
