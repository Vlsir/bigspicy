** Translated using xdm 2.6.0 on Nov_14_2022_16_05_25_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__pfet_g5v0d16v0 d g s b 
+ PARAMS: W=5.0 L=0.66 NF=1 AD=0 AS=0 PD=0 PS=0.0 M=1 NRD=0 NRS=0 SA=0.28 SB=1.19 SD=0 
+ MULT=1
.PARAM RDIFF='8.900000e+003*sky130_fd_pr__pfet_g5v0d16v0__rdiff_mult'
.PARAM RDIFF_TC1=2.500000e-003
.PARAM RDIFF_TC2=2.200000e-006
.PARAM SB_CADFIXEDVALUE_PVHV=1.19
* sd intentionally left out for sky130_fd_pr__pfet_g5v0d16v0 devices because poly-poly spacing not uniform in DE FET
Xmain1 d1 g s b sky130_fd_pr__pfet_g5v0d16v0__base 
+ PARAMS: W={w} L={l} NF={nf} AD=0 AS={as} PD=0 PS={ps} NRD={nrd} NRS={nrs} M={m} MULT={mult} 
+ SA={sa} SB={sb_cadfixedvalue_pvhv}
Rldd d d1 TC1='rdiff_tc1' TC2='rdiff_tc2' R='(1/w)*rdiff'
Dnw1 d b sky130_fd_pr__pfet_g5v0d16v0__parasitic__diode_pw2dn AREA='ad/2'
Dnw2 d1 b sky130_fd_pr__pfet_g5v0d16v0__parasitic__diode_pw2dn AREA='ad/2'
.ENDS sky130_fd_pr__pfet_g5v0d16v0
