** Translated using xdm 2.6.0 on Nov_14_2022_16_05_15_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 38
.PARAM 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__TOXE_MULT=1.052 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__OVERLAP_MULT=0.98026 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__AJUNCTION_MULT=1.1755 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__PJUNCTION_MULT=1.0477 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__RSHN_MULT=1.2 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__WINT_DIFF=3.2175e-8 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__DLC_DIFF=-1.5633e-8 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__DWC_DIFF=3.2175e-8 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__U0_DIFF_0=5.0533e-3 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__VSAT_DIFF_0=5.6551e+4 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__VTH0_DIFF_0=1.6480e-1 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__NFACTOR_DIFF_0=3.9755e-1 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__K2_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__UA_DIFF_0=0.0 SKY130_FD_PR__SPECIAL_NFET_PASS_LVT__UB_DIFF_0=0.0
*
* sky130_fd_pr__special_nfet_pass_lvt, Bin 000, W = 0.30, L = 0.15
* -------------------------------------
.INCLUDE sky130_fd_pr__special_nfet_pass_lvt.pm3.spice









