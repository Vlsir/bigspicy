** Translated using xdm 2.6.0 on Nov_14_2022_16_05_18_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
.INCLUDE sky130_fd_pr__nfet_01v8__ff.pm3.spice
.INCLUDE sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.INCLUDE sky130_fd_pr__nfet_01v8_lvt__ff.corner.spice
.INCLUDE sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.INCLUDE sky130_fd_pr__pfet_01v8__ff.corner.spice
.INCLUDE sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.INCLUDE sky130_fd_pr__nfet_03v3_nvt__ff.corner.spice
.INCLUDE sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
.INCLUDE sky130_fd_pr__nfet_05v0_nvt__ff.corner.spice
.INCLUDE sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.INCLUDE sky130_fd_pr__esd_nfet_01v8__ff.corner.spice
.INCLUDE sky130_fd_pr__pfet_01v8_lvt__ff.corner.spice
.INCLUDE sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.INCLUDE sky130_fd_pr__pfet_01v8_hvt__ff.pm3.spice
.INCLUDE sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.INCLUDE sky130_fd_pr__esd_pfet_g5v0d10v5__ff.corner.spice
.INCLUDE sky130_fd_pr__pfet_g5v0d10v5__ff.corner.spice
.INCLUDE sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.INCLUDE sky130_fd_pr__pfet_g5v0d16v0__ff.corner.spice
.INCLUDE sky130_fd_pr__nfet_g5v0d10v5__ff.corner.spice
.INCLUDE sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.INCLUDE sky130_fd_pr__nfet_g5v0d16v0__ff_discrete.corner.spice
.INCLUDE sky130_fd_pr__esd_nfet_g5v0d10v5__ff.corner.spice
.INCLUDE nonfet.spice
.INCLUDE sky130_fd_pr__pfet_20v0__fs_discrete.corner.spice
.INCLUDE sky130_fd_pr__nfet_20v0__sf_discrete.corner.spice
.INCLUDE sky130_fd_pr__nfet_20v0_nvt__sf_discrete.corner.spice
.INCLUDE all.spice
.INCLUDE rf.spice
