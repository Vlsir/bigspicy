** Translated using xdm 2.6.0 on Nov_14_2022_16_05_31_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 05
.PARAM 
+ SKY130_FD_PR__NFET_G5V0D16V0__TOXE_MULT=0.94 SKY130_FD_PR__NFET_G5V0D16V0__TOXP_MULT=1.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__OVERLAP_MULT=0.10246 SKY130_FD_PR__NFET_G5V0D16V0__AJUNCTION_MULT=8.1753e-1 
+ SKY130_FD_PR__NFET_G5V0D16V0__PJUNCTION_MULT=7.7786e-1 SKY130_FD_PR__NFET_G5V0D16V0__RDIFF_MULT=6.4330e-1 
+ SKY130_FD_PR__NFET_G5V0D16V0__LINT_DIFF=1.7325e-8 SKY130_FD_PR__NFET_G5V0D16V0__DLC_DIFF=1.7325e-8 
+ SKY130_FD_PR__NFET_G5V0D16V0__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__NFET_G5V0D16V0__DWC_DIFF=-3.2175e-8 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_0=-1.3425e-1 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_0=2.2191e-2 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_0=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_1=-0.14054 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_1=0.015572 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_1=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_2=-0.13714 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_2=0.016601 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_2=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_3=-0.097324 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_3=0.004226 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_3=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__VTH0_DIFF_4=-0.090898 SKY130_FD_PR__NFET_G5V0D16V0__U0_DIFF_4=0.0020803 
+ SKY130_FD_PR__NFET_G5V0D16V0__K2_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VSAT_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UA_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__UB_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__NFACTOR_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KT2_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__UTE_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__ETA0_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__DSUB_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__AGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_G5V0D16V0__CGIDL_DIFF_4=0.0 SKY130_FD_PR__NFET_G5V0D16V0__KETA_DIFF_4=0.0
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 000, W = 20.0, L = 0.7
* --------------------------------
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 001, W = 5.0, L = 0.7
* --------------------------------
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 002, W = 50.0, L = 0.7
* --------------------------------
*
















* sky130_fd_pr__nfet_g5v0d16v0, Bin 003, W = 20.0, L = 2.2
* --------------------------------
*






















* sky130_fd_pr__nfet_g5v0d16v0, Bin 004, W = 20.0, L = 2.2
* --------------------------------
.INCLUDE sky130_fd_pr__nfet_g5v0d16v0__subcircuit.pm3.spice






















.INCLUDE sky130_fd_pr__nfet_g5v0d16v0.pm3.spice
