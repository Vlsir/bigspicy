** Translated using xdm 2.6.0 on Nov_14_2022_16_05_14_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 9
.PARAM 
+ SKY130_FD_PR__NFET_03V3_NVT__TOXE_MULT=1.0365 SKY130_FD_PR__NFET_03V3_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_03V3_NVT__OVERLAP_MULT=1.1614 SKY130_FD_PR__NFET_03V3_NVT__AJUNCTION_MULT=1.2643 
+ SKY130_FD_PR__NFET_03V3_NVT__PJUNCTION_MULT=1.1856 SKY130_FD_PR__NFET_03V3_NVT__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__WINT_DIFF=2.252e-8 SKY130_FD_PR__NFET_03V3_NVT__DLC_DIFF=-3.0000e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__DWC_DIFF=2.252e-8 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_0=0.056603 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_0=0.018609 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_0=-1.6806 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_0=0.011726 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_0=-0.003049 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_0=-6511.3 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_0=1.7149e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_0=-2.5717e-11 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_1=-4.8514e-12 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_1=0.048996 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_1=0.018393 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_1=-1.4856 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_1=0.019978 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_1=-0.0035858 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_1=-3705.6 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_1=3.9763e-19 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_2=3.9604e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_2=8.898e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_2=0.0099926 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_2=-0.42593 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_2=0.040995 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_2=0.006932 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_2=507.3 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_3=-4.3506e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_3=-5.8077e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_3=0.060669 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_3=0.018737 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_3=-1.7015 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_3=0.0082446 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_3=-0.0029241 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_3=-5671.4 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_4=3.1881e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_4=-1.0615e-10 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_4=0.030291 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_4=0.010253 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_4=-1.1697 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_4=0.043806 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_4=-0.0071731 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_4=-13214.0 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_5=0.0012881 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_5=-11299.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_5=4.4342e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_5=-4.5129e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_5=0.019094 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_5=-1.6081 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_5=0.08882 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_6=-0.67715 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_6=0.048142 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_6=0.00057016 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_6=-5077.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_6=2.8143e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_6=1.972e-10 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_6=0.017779 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_7=0.05271 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_7=0.018319 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_7=-1.4409 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_7=0.023503 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_7=-0.0051263 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_7=-6539.7 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_7=1.5451e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_7=-1.5534e-10 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_8=0.012232 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_8=-0.3358 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_8=0.034016 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_8=0.0036844 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_8=-1219.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_8=3.1622e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_8=7.4928e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_8=0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
*














* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_03v3_nvt.pm3.spice




















