** Translated using xdm 2.6.0 on Nov_14_2022_16_05_32_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TOXE_MULT=1.06 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RSHP_MULT=1.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__OVERLAP_MULT=1.292 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AJUNCTION_MULT=1.0777e+0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PJUNCTION_MULT=1.0736e+0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__WINT_DIFF=3.2175e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__DLC_DIFF=-1.7325e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__DWC_DIFF=3.2175e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_0=8.3700e-3 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_0=2.6732e-3 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_0=9.4633e+4 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_0=-5.8555e-2 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_0=-4.2555e-1 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_0=1.9037e-10 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_0=1.0572e-18 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_0=-1.1583e-3 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_1=0.15309 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_1=0.015841 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_1=-0.0066616 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_1=22080.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_1=0.070909 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_1=-5.5136e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_1=0.51452 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_1=-3.0377e-18 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_2=5.4092e-2 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_2=1.0843e-2 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_2=2.4584e-4 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_2=-2.9721e-2 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_2=3.6720e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_2=6.4607e+4 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_2=3.7549e-1 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_2=1.9733e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_3=3.3063e-2 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_3=9.1109e-3 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_3=2.0202e-3 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_3=-5.2973e-2 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_3=7.2069e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_3=4.3170e+4 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_3=1.2833e-1 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_3=7.6394e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_4=0.022785 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_4=0.0088938 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_4=0.0020785 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_4='-0.06018-0.005' SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_4=5.9115e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_4=47898.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_4=-0.1672 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_4=9.8318e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_5=0.16248 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_5=0.016552 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_5=-0.0073777 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_5=0.078938 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_5=-5.267e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_5=28612.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_5=0.56919 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_5=-3.3626e-18 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_6=-3.936e-18 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_6=0.18617 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_6=0.016075 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_6=-0.0087419 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_6=0.11079 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_6=-4.0545e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_6=40444.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_6=0.47252 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_7=-2.7759e-18 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_7=0.14442 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_7=0.016523 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_7=-0.006295 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_7=0.059613 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_7=1.6811e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_7=21388.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_7=0.57083 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_7=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
*




* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
.INCLUDE sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice























