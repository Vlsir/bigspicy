** Translated using xdm 2.6.0 on Nov_14_2022_16_05_04_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PFET_01V8__TOXE_SLOPE=4.443e-03
.PARAM SKY130_FD_PR__PFET_01V8__TOXE_SLOPE1=6.443e-03
.PARAM SKY130_FD_PR__PFET_01V8__TOXE_SLOPE2=3.443e-03
.PARAM SKY130_FD_PR__PFET_01V8__LINT_SLOPE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE=0.1
.PARAM SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE1=0.1
.PARAM SKY130_FD_PR__PFET_01V8__NFACTOR_SLOPE2=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VOFF_SLOPE=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VOFF_SLOPE1=0.0
.PARAM SKY130_FD_PR__PFET_01V8__VOFF_SLOPE2=0.007
.PARAM SKY130_FD_PR__PFET_01V8__VTH0_SLOPE=5.856e-03
.PARAM SKY130_FD_PR__PFET_01V8__VTH0_SLOPE1=7.356e-03
.PARAM SKY130_FD_PR__PFET_01V8__VTH0_SLOPE2=4.356e-03
.PARAM SKY130_FD_PR__PFET_01V8__WINT_SLOPE=0
