** Translated using xdm 2.6.0 on Nov_14_2022_16_05_28_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.INCLUDE 
+ sky130_fd_pr__nfet_20v0_zvt__parasitic__diode_ps2dn__extended_drain.model.spice
.SUBCKT sky130_fd_pr__nfet_20v0_zvt d g s b 
+ PARAMS: W=60u L=2u M=1 T=30 AD=0 AS=0 PD=0 PS=0 NRD=2 NRS=2 MF=1 SA=0 SB=0
.PARAM 
+ RDRIFT_TNOM=4.73057453e+003 VGDEP_TNOM=0.020646 VTH_TNOM=7.000000e-001 VBDEP_TNOM=-5.260300e-001 
+ VTH2=0.5 HVVSAT_TNOM=1.236813882 AVSAT_TNOM=7.467500e-001 DELTAW=9.000000e-001 
+ HVNEL_N20ZVTVHV1=5.00 HVVBDEP=-2.490600e-002
.PARAM 
+ SKY130_FD_PR__NFET_20V0_ZVT__PGATEJUNCTION_MULT=1.7357 SKY130_FD_PR__NFET_20V0_ZVT__MJSWGATEJUNCTION_MULT=5.3981e-1 
+ SKY130_FD_PR__NFET_20V0_ZVT__PBSWGATEJUNCTION_MULT=3.4999e+0
.PARAM 
+ SKY130_FD_PR__NFET_20V0_ZVT__VGDEP_MULT=1 N20ZVTVHV1RES_VTH0_DIFF=0.0 SKY130_FD_PR__NFET_20V0_ZVT__VBDEP_MULT=1 
+ SKY130_FD_PR__NFET_20V0_ZVT__AVSAT_MULT=0.984
.PARAM 
+ W_N20ZVTVHV1=30.00 NRD_N20ZVTVHV1=2.0 NRS_N20ZVTVHV1=2.0 AD_N20ZVTVHV1=103.5 AS_N20ZVTVHV1=8.7 
+ PD_N20ZVTVHV1=41.75 PS_N20ZVTVHV1=60.58 DELVTO_N20ZVTVHV1=0.0
.PARAM TC1_VGDEP=0






.PARAM TC1_VTH=0
.PARAM TC1_VBDEP=0
.PARAM TC1_HVVSAT_N20ZVTVHV1=0.0061411164700097
.PARAM TC2_RDRIFT_N20ZVTVHV1=5.0768e-005
.PARAM TC2_VGDEP=0
.PARAM TC2_VTH=0
.PARAM TC2_VBDEP=0
.PARAM TC2_HVVSAT_N20ZVTVHV1=3.61396725197052E-05
.PARAM TC2_AVSAT_N20ZVTVHV1=3.0122688512968E-06
.PARAM TC1_RDRIFT_N20ZVTVHV1=0.012359
.PARAM TC1_AVSAT_N20ZVTVHV1=-7.4563e-04
.PARAM 
+ RDRIFT='rdrift_tnom*((w_n20zvtvhv1-deltaw)/w_n20zvtvhv1)*(1+tc1_rdrift_n20zvtvhv1*(temp-30)+tc2_rdrift_n20zvtvhv1*(temp-30)*(temp-30))*sky130_fd_pr__nfet_20v0_zvt__rdrift_mult' 
+ VGDEP='vgdep_tnom*(1+tc1_vgdep*(temp-30)+tc2_vgdep*(temp-30)*(temp-30))*sky130_fd_pr__nfet_20v0_zvt__vgdep_mult' 
+ VTH='vth_tnom*(1+tc1_vth*(temp-30)+tc2_vth*(temp-30)*(temp-30))+n20zvtvhv1res_vth0_diff' 
+ VBDEP='vbdep_tnom*(1+tc1_vbdep*(temp-30)+tc2_vbdep*(temp-30)*(temp-30))*sky130_fd_pr__nfet_20v0_zvt__vbdep_mult' 
+ HVVSAT='hvvsat_tnom*(1+tc1_hvvsat_n20zvtvhv1*(temp-30)+tc2_hvvsat_n20zvtvhv1*(temp-30)*(temp-30))*sky130_fd_pr__nfet_20v0_zvt__hvvsat_mult' 
+ AVSAT='avsat_tnom*(1+tc1_avsat_n20zvtvhv1*(temp-30)+tc2_avsat_n20zvtvhv1*(temp-30)*(temp-30))*sky130_fd_pr__nfet_20v0_zvt__avsat_mult'
M1 d1 g s b sky130_fd_pr__nfet_20v0_zvt__base 
+ M={m} AD=0 AS=0 L={hvnel_n20zvtvhv1} NRD={nrd_n20zvtvhv1} NRS={nrs_n20zvtvhv1} 
+ PD=0 PS=0 W={w_n20zvtvhv1}
* rldd d d1 r='abs((1/w_n20zvtvhv1)*(rdrift/(1+vgdep*(v(g,s)-vth-vbdep*v(b,s))))*(1+pwr((abs(v(d,s)+vth2-min(v(d1,s),60))/(hvvsat*(1+hvvbdep*v(b,s)))),avsat)))' tc1 = 0 tc2 = 0 m = {m}; HSpice Parser Retained (as a comment). Continuing.
DNDrain1 b d sky130_fd_pr__nfet_20v0_zvt__parasitic__diode_ps2dn__extended_drain 
+ AREA='0.5*ad_n20zvtvhv1'
DNDrain2 b d1 
+ sky130_fd_pr__nfet_20v0_zvt__parasitic__diode_ps2dn__extended_drain 
+ AREA='0.5*ad_n20zvtvhv1'
DNSrc b s sky130_fd_pr__diode_pw2nd_05v5 AREA={as_n20zvtvhv1}
* DC IV MOS Parameters
* BSIM4 - Model Selectors




















* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters













.ENDS sky130_fd_pr__nfet_20v0_zvt





















*.END
