** Translated using xdm 2.6.0 on Nov_14_2022_16_05_14_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__TOXE_MULT=1.0365 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__OVERLAP_MULT=9.6320e-1 SKY130_FD_PR__RF_NFET_01V8_LVT_B__AJUNCTION_MULT=1.1229e+0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__PJUNCTION_MULT=1.0009e+0 SKY130_FD_PR__RF_NFET_01V8_LVT_B__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__WINT_DIFF=2.252e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__DLC_DIFF=-1.1228e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__XGW_DIFF=4.504e-8 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT_P42=1.1125 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT_P42=1.245 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT_P42=1.245 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT=1.1125 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT=1.245 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT=1.245 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RS_MULT=1.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_0=0.035472 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_0=-0.0035791 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_0=11669.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_0=-0.023208 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_1=-0.015447 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_1=0.031659 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_1=-0.0022517 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_1=16627.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_2=-0.00027242 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_2=0.006014 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_2=-0.0024036 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_2=7476.5 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_3=-0.025698 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_3=0.022412 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_3=-0.0067063 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_3=14950.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_4=-0.018667 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_4=0.0074967 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_4=-0.0031604 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_4=14641.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_5=-0.0050153 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_5=0.005408 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_5=-0.0036655 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_5=14592.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_6=-0.031185 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_6=0.019026 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_6=-0.0097006 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_6=9042.7 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_7=-0.018406 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_7=0.005177 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_7=-0.0054184 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_7=13962.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_8=-0.0045172 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_8=0.0026993 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_8=-0.0049523 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_8=16409.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_0=-0.022384 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_0=0.032174 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_0=-0.0088162 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_0=18475.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_1=-0.015672 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_1=0.024627 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_1=-0.0052084 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_1=17204.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_2=-0.0053553 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_2=0.00058529 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_2=-0.0047533 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_2=14144.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_3=-0.026679 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_3=0.025797 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_3=-0.0070348 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_3=14175.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_4=-0.007826 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_4=18436.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_4=-0.019062 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_4=0.0093971 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_5=-0.0078718 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_5=-0.0066522 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_5=26781.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_5=-0.0060231 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_6=-0.03107 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_6=0.017691 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_6=-0.0077169 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_6=12148.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_7=-0.019933 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_7=0.0024544 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_7=-0.0097882 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_7=13883.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_8=-0.0057624 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_8=-0.0093065 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_8=39684.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_8=-0.014919 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_8=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice















