** Translated using xdm 2.6.0 on Nov_14_2022_16_05_16_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__TOXE_MULT=1.052 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__OVERLAP_MULT=9.8026e-1 SKY130_FD_PR__RF_NFET_01V8_LVT_B__AJUNCTION_MULT=1.1755e+0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__PJUNCTION_MULT=1.0477e+0 SKY130_FD_PR__RF_NFET_01V8_LVT_B__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__WINT_DIFF=3.2175e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__DLC_DIFF=-1.5633e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__XGW_DIFF=6.4250e-8 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT_P42=1.15 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT_P42=1.35 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT_P42=1.35 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT=1.15 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT=1.35 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT=1.35 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RS_MULT=1.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_0=0.053368 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_0=-0.0019719 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_0=26569.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_0=-0.024863 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_1=-0.017808 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_1=0.047766 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_1=-0.00047355 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_1=30213.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_2=0.00040478 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_2=0.015345 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_2=-0.001204 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_2=18070.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_3=-0.029988 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_3=0.037878 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_3=-0.0051828 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_3=28757.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_4=-0.022408 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_4=0.020083 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_4=-0.0014964 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_4=25513.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_5=-0.0063582 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_5=0.012 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_5=-0.0026836 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_5=24731.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_6=-0.034961 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_6=0.032444 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_6=-0.0082913 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_6=19960.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_7=-0.021804 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_7=0.01554 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_7=-0.0040633 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_7=23539.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_8=-0.0057548 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_8=0.0080085 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_8=-0.0040879 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_8=26010.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_0=-0.023869 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_0=0.050138 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_0=-0.0074552 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_0=34785.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_1=-0.017943 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_1=0.040645 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_1=-0.0035828 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_1=30760.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_2=-0.0065733 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_2=0.009983 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_2=-0.0036611 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_2=24896.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_3=-0.030893 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_3=0.041356 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_3=-0.0055014 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_3=28064.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_4=-0.0064683 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_4=30230.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_4=-0.022603 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_4=0.021578 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_5=-0.0014353 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_5=-0.0058089 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_5=37969.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_5=-0.0073485 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_6=-0.035237 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_6=0.031623 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_6=-0.0062253 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_6=24780.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_7=-0.02312 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_7=0.012306 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_7=-0.0086402 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_7=24437.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_8=-0.0069151 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_8=-0.0086411 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_8=52788.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_8=-0.0097748 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_8=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice















