** Translated using xdm 2.6.0 on Nov_14_2022_16_05_18_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 9
.PARAM 
+ SKY130_FD_PR__NFET_03V3_NVT__TOXE_MULT=1.052 SKY130_FD_PR__NFET_03V3_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_03V3_NVT__OVERLAP_MULT=1.37 SKY130_FD_PR__NFET_03V3_NVT__AJUNCTION_MULT=1.3878 
+ SKY130_FD_PR__NFET_03V3_NVT__PJUNCTION_MULT=1.2464 SKY130_FD_PR__NFET_03V3_NVT__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__WINT_DIFF=3.2175e-8 SKY130_FD_PR__NFET_03V3_NVT__DLC_DIFF=-3.0000e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__DWC_DIFF=3.2175e-8 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_0=0.070007 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_0=0.025405 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_0=-1.8 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_0=0.01866 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_0=-0.0034806 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_0=-4720.5 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_0=-1.0e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_0=1.1794e-11 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_1=7.2867e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_1=0.061113 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_1=0.022045 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_1=-1.5295 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_1=0.030601 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_1=-0.00236 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_1=937.82 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_1=-7.7567e-19 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_2=4.3331e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_2=8.8389e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_2=0.0117 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_2=-0.4369 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_2=0.057242 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_2=0.011419 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_2=5633.8 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_3=-2.5164e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_3=9.4843e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_3=0.077321 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_3=0.024946 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_3=-1.8358 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_3=0.012417 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_3=-0.0043072 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_3=-3550.1 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_4=4.2773e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_4=1.029e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_4=0.017434 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_4=0.0092175 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_4=-1.2004 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_4=0.076144 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_4=0.0014096 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_4=-4990.9 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_5=0.0070104 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_5=-3975.1 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_5=4.2056e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_5=1.6413e-10 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_5=0.021544 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_5=-1.6491 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_5=0.10543 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_6=-0.70119 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_6=0.059414 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_6=0.0049892 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_6=2172.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_6=2.8836e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_6=2.4441e-10 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_6=0.020119 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_7=0.069322 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_7=0.021677 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_7=-1.4753 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_7=0.028831 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_7=-0.0053542 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_7=-1407.8 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_7=-4.6026e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_7=-2.6093e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_8=0.013898 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_8=-0.33169 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_8=0.050109 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_8=0.0080728 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_8=4767.8 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_8=3.6297e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_8=-2.7576e-13 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_8=0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
*














* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_03v3_nvt.pm3.spice




















