** Translated using xdm 2.6.0 on Nov_14_2022_16_05_17_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TOXE_MULT=1.06 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RSHN_MULT=1.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__OVERLAP_MULT=1.0412 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AJUNCTION_MULT=1.1726e+0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PJUNCTION_MULT=1.2510e+0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__LINT_DIFF=-1.7325e-8 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__WINT_DIFF=3.2175e-8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__DLC_DIFF=-1.7325e-8 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__DWC_DIFF=3.2175e-8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_0=0.32023 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_0=0.020037 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_0=0.002635 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_0=0.029648 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_0=4367.2 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_0=1.509e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_0=6.7217e-13 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_1=0.30154 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_1=0.019119 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_1=0.0043558 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_1=0.030739 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_1=4689.7 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_1=1.6267e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_1=-1.2957e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_2=0.29898 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_2=0.019424 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_2=0.0025388 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_2=0.030149 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_2=5961.9 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_2=1.6089e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_2=-3.8247e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_3=6.5182e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_3=0.30517 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_3=0.01879 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_3=0.0023371 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_3=0.028108 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_3=6027.6 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_3=1.5974e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_4=1.5634e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_4=4.9713e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_4=0.30409 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_4=0.021181 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_4=0.0027289 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_4=0.027395 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_4=5017.5 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_5=-1.2342e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_5=5.7749e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_5=0.35342 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_5=0.10245 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_5=0.15639 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_5=0.042547 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_5=-0.0070149 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_5=0.014756 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_6=1.9501e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_6=3.7828e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_6=0.30885 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_6=0.019873 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_6=0.0030646 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_6=0.026727 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_6=7814.9 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_7=9619.4 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_7=2.3893e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_7=1.2122e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_7=0.27258 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_7=0.020512 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_7=0.0028097 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_7=0.026182 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_8=-0.0090729 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_8=-0.0044111 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_8=-1.0249e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_8=5.8119e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_8=0.33378 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_8=0.14336 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_8=0.21714 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_8=0.007425 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_9=0.0079697 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_9=0.0052236 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_9=0.016479 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_9=6132.2 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_9=2.7471e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_9=2.2591e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_9=0.2845 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_10=4.3397e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_10=2578.9 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_10=8.2269e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_10=0.0087889 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_10=0.31183 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_10=0.0011957 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_10=0.028866 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
*
















* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
.INCLUDE sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice























