** Translated using xdm 2.6.0 on Nov_14_2022_16_05_03_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TOXE_MULT=1.042 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RSHN_MULT=1.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__OVERLAP_MULT=0.99758 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AJUNCTION_MULT=1.1193e+0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PJUNCTION_MULT=1.1801e+0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__WINT_DIFF=2.252e-8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__DLC_DIFF=-1.21275e-8 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__DWC_DIFF=2.252e-8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_0=0.30329 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_0=0.01726 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_0=0.00068868 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_0=0.024431 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_0=1583.3 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_0=1.32e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_0=1.6741e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_1=0.28901 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_1=0.01659 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_1=0.0023767 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_1=0.025579 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_1=1895.9 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_1=1.438e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_1=2.8248e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_2=0.28823 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_2=0.016801 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_2=0.00060123 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_2=0.024939 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_2=3195.6 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_2=1.4202e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_2=1.0136e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_3=1.3648e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_3=0.29555 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_3=0.016145 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_3=0.00028215 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_3=0.023983 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_3=3192.2 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_3=1.3881e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_4=1.3703e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_4=1.7829e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_4=0.2895 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_4=0.017958 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_4=0.00077795 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_4=0.022447 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_4=2279.7 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_5=-2.1985e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_5=6.9289e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_5=0.33754 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_5=0.049359 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_5=0.071277 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_5=0.043943 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_5=-0.0080434 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_5=0.013646 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_6=1.7407e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_6=1.9509e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_6=0.29323 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_6=0.017035 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_6=0.0011167 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_6=0.021986 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_6=4980.3 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_7=6726.2 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_7=2.17e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_7=1.9011e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_7=0.25951 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_7=0.017543 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_7=0.00080633 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_7=0.021766 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_8=-0.010132 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_8=-0.0032051 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_8=-2.1641e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_8=6.8574e-11 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_8=0.31944 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_8=0.10492 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_8=0.15983 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_8=0.00845 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_9=0.0060854 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_9=0.0032612 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_9=0.012301 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_9=3335.1 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_9=2.5113e-18 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_9=1.4426e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_9=0.27036 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_10=1.0694e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_10=-198.96 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_10=7.208e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_10=0.0071747 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_10=0.31463 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_10=-0.00052628 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_10=0.024124 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
*
















* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
.INCLUDE sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice























