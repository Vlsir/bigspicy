** Translated using xdm 2.6.0 on Nov_14_2022_16_05_34_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* SKY130 Spice File.
* Typical Varactor Parameters
.PARAM 
+ CNWVC_TOX='41.6503*1.024' CNWVC_CDEPMULT=1 CNWVC_CINTMULT=1 CNWVC_VT1=0.3333 CNWVC_VT2=0.2380952 
+ CNWVC_VTR=0.16 CNWVC_DWC=0.0 CNWVC_DLC=0.0 CNWVC_DLD=0.0 CNWVC2_TOX='41.7642*1.017' 
+ CNWVC2_CDEPMULT=1 CNWVC2_CINTMULT=1 CNWVC2_VT1=0.2 CNWVC2_VT2=0.33 CNWVC2_VTR=0.14 
+ CNWVC2_DWC=0.0 CNWVC2_DLC=0.0 CNWVC2_DLD=0.0
* sky130_fd_pr__model__parasitic__diode_ps2nw Parameters














* .param  sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 9.8286e-01    ; Units: farad/meter^2   sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 9.8954e-01    ; Units: farad/meter^2   sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult = 9.8580e-01  ; Units: farad/meter   sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 1.0116e+0   ; Units: farad/meter   sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 9.8200e-01      ; Units: farad/meter   sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult = 9.6304e-01       ; Units: farad/meter   sky130_fd_pr__nfet_01v8__ajunction_mult = 9.9543e-1   sky130_fd_pr__nfet_01v8__pjunction_mult = 1.0204e+0   sky130_fd_pr__pfet_01v8_hvt__ajunction_mult = 9.8366e-1   sky130_fd_pr__pfet_01v8_hvt__pjunction_mult = 1.0286e+0   dkispp=9.2840e-01 dkbfpp=9.5154e-01 dknfpp=1.000   dkispp5x=1.0046e+00 dkbfpp5x=1.1288e+00 dknfpp5x=1.0009e+00 dkisepp5x=0.745   cvpp2_nhvnative10x4_cor=1.00   cvpp2_nhvnative10x4_sub=4.82e-15   cvpp2_phv5x4_cor=1.00   cvpp2_phv5x4_sub=4.82e-15; HSpice Parser Retained (as a comment). Continuing.
* sky130_fd_pr__model__parasitic__diode_ps2dn Parameters


* sky130_fd_pr__model__parasitic__diode_pw2dn Parameters


* sky130_fd_pr__diode_pw2nd_05v5  Parameters


* sky130_fd_pr__diode_pd2nw_05v5_hvt  Parameters


