** Translated using xdm 2.6.0 on Nov_14_2022_16_05_31_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 9
.PARAM 
+ SKY130_FD_PR__NFET_03V3_NVT__TOXE_MULT=0.948 SKY130_FD_PR__NFET_03V3_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_03V3_NVT__OVERLAP_MULT=0.40927 SKY130_FD_PR__NFET_03V3_NVT__AJUNCTION_MULT=0.56418 
+ SKY130_FD_PR__NFET_03V3_NVT__PJUNCTION_MULT=0.84099 SKY130_FD_PR__NFET_03V3_NVT__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__NFET_03V3_NVT__DLC_DIFF=3.0000e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__DWC_DIFF=-3.2175e-8 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_0=-0.0010542 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_0=-0.026492 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_0=-1.0339 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_0=-0.047264 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_0=0.00016819 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_0=-3949.2 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_0=4.2013e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_0=5.9282e-11 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_1=8.318e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_1=-0.020875 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_1=-0.0056301 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_1=-1.707 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_1=-0.060897 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_1=-0.0028636 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_1=-14012.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_1=4.2893e-19 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_2=1.0603e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_2=4.1221e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_2=-0.00080074 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_2=-0.47778 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_2=-0.050539 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_2=-0.00039963 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_2=-12436.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_3=7.9696e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_3=5.7902e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_3=-0.0026756 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_3=-0.023644 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_3=-0.95532 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_3=-0.048464 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_3=0.0011558 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_3=-6147.9 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_4=1.7046e-19 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_4=3.9478e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_4=0.032977 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_4=0.0069451 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_4=-1.6941 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_4=-0.083671 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_4=-0.0011543 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_4=-12626.0 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_5=0.0089834 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_5=-11481.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_5=1.7135e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_5=4.1927e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_5=0.0029293 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_5=-1.5761 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_5=-0.0016017 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_6=-0.73851 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_6=-0.014966 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_6=0.0066129 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_6=-9425.6 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_6=1.5395e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_6=6.8955e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_6=0.0030242 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_7=-0.0078507 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_7=-0.0030712 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_7=-1.5397 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_7=-0.053605 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_7=-0.000432 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_7=-14226.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_7=1.2313e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_7=6.9284e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_8=0.0019101 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_8=-0.52333 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_8=-0.057025 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_8=0.00086474 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_8=-12780.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_8=1.3078e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_8=4.5353e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_8=0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
*














* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_03v3_nvt.pm3.spice




















