** Translated using xdm 2.6.0 on Nov_14_2022_16_05_06_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PFET_01V8_HVT__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_HVT__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_HVT__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_HVT__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__pfet_01v8_hvt d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__pfet_01v8_hvt d g s b sky130_fd_pr__pfet_01v8_hvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.095122+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43657182   k2 = 0.038826066   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.16832488+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5988376+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.009347598   ua = -5.257697e-11   ub = 7.671173e-20   uc = -7.7670696e-11   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 200000.0   a0 = 1.597986   ags = 0.2656338   a1 = 0.0   a2 = 1.0   b0 = 0.0   b1 = 0.0   keta = -0.013169082   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.075489662   pdiblc1 = 0.39   pdiblc2 = 0.0036275994   pdiblcb = -9.5744039e-5   drout = 0.56   pscbe1 = 746475130.0   pscbe2 = 9.5049925e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.7923891   agidl = 1.0e-10   bgidl = 1154444600.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.44169   kt2 = -0.037961   at = 0.0   ute = -0.30066   ua1 = 2.2116e-9   ub1 = -7.9359e-19   uc1 = 1.1985e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.095122+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43657182   k2 = 0.038826066   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.16832488+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.5988376+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.009347598   ua = -5.257697e-11   ub = 7.671173e-20   uc = -7.7670696e-11   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 200000.0   a0 = 1.597986   ags = 0.2656338   a1 = 0.0   a2 = 1.0   b0 = 0.0   b1 = 0.0   keta = -0.013169082   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.075489662   pdiblc1 = 0.39   pdiblc2 = 0.0036275994   pdiblcb = -9.5744039e-5   drout = 0.56   pscbe1 = 746475130.0   pscbe2 = 9.5049925e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.7923891   agidl = 1.0e-10   bgidl = 1154444600.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.44169   kt2 = -0.037961   at = 0.0   ute = -0.30066   ua1 = 2.2116e-9   ub1 = -7.9359e-19   uc1 = 1.1985e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.094651495e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.786514799e-09 wvth0 = -4.702045241e-08 pvth0 = 3.784100214e-13   k1 = 4.360523215e-01 lk1 = 4.180806759e-09 wk1 = 5.191671912e-08 pk1 = -4.178140742e-13   k2 = 3.905734125e-02 lk2 = -1.861251206e-09 wk2 = -2.311277742e-08 pk2 = 1.860064323e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.682664013e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.706235798e-10 wvoff = -5.844142915e-09 pvoff = 4.703234725e-14   nfactor = {1.594203349e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.729540931e-08 wnfactor = 4.631295827e-07 pnfactor = -3.727162678e-12   eta0 = 0.08   etab = -0.07   u0 = 9.359080907e-03 lu0 = -9.241185555e-11 wu0 = -1.147558504e-09 pu0 = 9.235292636e-15   ua = -4.920615129e-11 lua = -2.712759058e-17 wua = -3.368669211e-16 pua = 2.711029186e-21   ub = 7.263134604e-20 lub = 3.283801204e-26 wub = 4.077781983e-25 pub = -3.281707190e-30   uc = -7.712327301e-11 luc = -4.405537080e-18 wuc = -5.470739127e-17 puc = 4.402727758e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.943936016e+05 lvsat = 4.511903282e-02 wvsat = 5.602823304e-01 pvsat = -4.509026131e-6   a0 = 1.618382908e+00 la0 = -1.641497290e-07 wa0 = -2.038390164e-06 pa0 = 1.640450540e-11   ags = 2.847666745e-01 lags = -1.539770693e-07 wags = -1.912067388e-06 pags = 1.538788812e-11   a1 = 0.0   a2 = 9.848959663e-01 la2 = 1.214733870e-07 wa2 = 1.508440853e-06 pa2 = -1.213959259e-11   b0 = 0.0   b1 = 0.0   keta = -1.635496691e-02 lketa = 2.563928496e-08 wketa = 3.183853339e-07 pketa = -2.562293530e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.175530136e-01 lpclm = -3.385163897e-07 wpclm = -4.203652868e-06 ppclm = 3.383005246e-11   pdiblc1 = 0.39   pdiblc2 = 3.389891695e-03 lpdiblc2 = 1.913018123e-09 wpdiblc2 = 2.375561232e-08 ppdiblc2 = -1.911798230e-13   pdiblcb = -1.467140768e-04 lpdiblcb = 4.101953961e-10 wpdiblcb = 5.093753525e-09 ppdiblcb = -4.099338227e-14   drout = 0.56   pscbe1 = 7.505148629e+08 lpscbe1 = -3.251086178e+01 wpscbe1 = -4.037156886e+02 ppscbe1 = 3.249013026e-3   pscbe2 = 9.463149641e-09 lpscbe2 = 3.367419162e-16 wpscbe2 = 4.181617684e-15 ppscbe2 = -3.365271826e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.831940178e+00 lbeta0 = -3.182981755e-07 wbeta0 = -3.952585692e-06 pbeta0 = 3.180952032e-11   agidl = 1.034218799e-10 lagidl = -2.753851915e-17 wagidl = -3.419697791e-16 pagidl = 2.752095839e-21   bgidl = 1.142788057e+09 lbgidl = 9.380923379e+01 wbgidl = 1.164910966e+03 pbgidl = -9.374941352e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.425028544e-01 lkt1 = 6.541668973e-09 wkt1 = 8.123360161e-08 pkt1 = -6.537497482e-13   kt2 = -3.814100535e-02 lkt2 = 1.448642572e-09 wkt2 = 1.798905662e-08 pkt2 = -1.447718802e-13   at = 1.981266456e+04 lat = -1.594478665e-01 wat = -1.980003042e+00 pat = 1.593461898e-5   ute = -3.004781078e-01 lute = -1.463827505e-09 wute = -1.817762116e-08 pute = 1.462894051e-13   ua1 = 2.227208011e-09 lua1 = -1.256097626e-16 wua1 = -1.559805832e-15 pua1 = 1.255296638e-20   ub1 = -8.067398249e-19 lub1 = 1.058268324e-25 wub1 = 1.314143956e-24 pub1 = -1.057593488e-29   uc1 = 1.211383402e-10 luc1 = -1.036827199e-17 wuc1 = -1.287518644e-16 puc1 = 1.036166035e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.101852341e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.536088631e-08 wvth0 = 3.472044050e-08 pvth0 = 4.754127859e-14   k1 = 4.496343333e-01 lk1 = -5.079612074e-08 wk1 = -6.011106403e-07 pk1 = 2.225493746e-12   k2 = 3.333508785e-02 lk2 = 2.130114307e-08 wk2 = 2.351972778e-07 pk2 = -8.595745513e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 5.440048812e-01 ldsub = 6.474464217e-08 wdsub = 1.598491907e-06 pdsub = -6.470335581e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.687524048e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.496609471e-09 wvoff = -3.655704093e-08 pvoff = 1.713512480e-13   nfactor = {1.695254432e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.717366399e-07 wnfactor = -3.352669920e-06 pnfactor = 1.171833515e-11   eta0 = 7.392900281e-02 leta0 = 2.457403065e-08 weta0 = 6.067125837e-07 peta0 = -2.455836029e-12   etab = -6.469265025e-02 letab = -2.148295762e-08 wetab = -5.303965355e-07 petab = 2.146925836e-12   u0 = 9.039325974e-03 lu0 = 1.201884170e-09 wu0 = 1.523964440e-08 pu0 = -5.709641761e-14   ua = -1.370214031e-10 lua = 3.283287903e-16 wua = 3.869086096e-15 pua = -1.431372229e-20   ub = 1.586658892e-19 lub = -3.154104611e-25 wub = -2.658227606e-24 pub = 9.128794454e-30   uc = -8.637304797e-11 luc = 3.303547075e-17 wuc = 1.275139958e-16 puc = -2.973183991e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.820211026e+05 lvsat = -3.095773749e-01 wvsat = -5.960304494e-01 pvsat = 1.714678307e-7   a0 = 1.280891365e+00 la0 = 1.201940104e-06 wa0 = 4.036225980e-06 pa0 = -8.184173961e-12   ags = -1.911761452e-02 lags = 1.076078159e-06 wags = 2.517674546e-06 pags = -2.542710533e-12   a1 = 0.0   a2 = 1.234945329e+00 la2 = -8.906701701e-07 wa2 = -3.016881706e-06 pa2 = 6.177894935e-12   b0 = 0.0   b1 = 0.0   keta = 3.624649252e-02 lketa = -1.872795875e-07 wketa = -6.191571299e-07 pketa = 1.232667416e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.810850624e-01 lpclm = 2.489413349e-06 wpclm = 8.588403566e-06 ppclm = -1.794931377e-11   pdiblc1 = 0.39   pdiblc2 = 7.309897997e-03 lpdiblc2 = -1.395428538e-08 wpdiblc2 = -4.572389188e-08 ppdiblc2 = 9.005757717e-14   pdiblcb = 6.389588179e-04 lpdiblcb = -2.770031705e-09 wpdiblcb = -4.321034876e-09 ppdiblcb = -2.884437151e-15   drout = 0.56   pscbe1 = 6.835922188e+08 lpscbe1 = 2.383769442e+02 wpscbe1 = 8.074313771e+02 ppscbe1 = -1.653437788e-3   pscbe2 = 1.013508658e-08 lpscbe2 = -2.383107626e-15 wpscbe2 = -6.240959330e-15 ppscbe2 = 8.535528414e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.327591634e+00 lbeta0 = 1.723191250e-06 wbeta0 = -7.171089136e-06 pbeta0 = 4.483729809e-11   agidl = 4.367544253e-11 lagidl = 2.143016162e-16 wagidl = 9.896657686e-16 pagidl = -2.638065240e-21   bgidl = 1.335891581e+09 lbgidl = -6.878303823e+02 wbgidl = -2.329821933e+03 pbgidl = 4.770951108e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.273730351e-01 lkt1 = -5.470043506e-08 wkt1 = -3.287598724e-07 pkt1 = 1.005811586e-12   kt2 = -3.541468677e-02 lkt2 = -9.586881614e-09 wkt2 = -1.042750029e-08 pkt2 = -2.974805152e-14   at = -3.215109905e+05 lat = 1.222153492e+00 wat = 5.269665788e+00 pat = -1.341040927e-5   ute = -2.934389274e-01 lute = -2.995684595e-08 wute = -9.682463222e-07 pute = 3.991953742e-12   ua1 = 1.924108124e-09 lua1 = 1.101270385e-15 wua1 = 7.570363599e-15 pua1 = -2.440390519e-20   ub1 = -5.635972638e-19 lub1 = -8.783595479e-25 wub1 = -5.156791224e-24 pub1 = 1.561695477e-29   uc1 = 8.381738267e-11 luc1 = 1.406985669e-16 wuc1 = 1.854302565e-15 puc1 = -6.990792106e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.090247229e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.596228745e-09 wvth0 = 1.358362197e-07 pvth0 = -1.595210862e-13   k1 = 4.209018192e-01 lk1 = 8.041603203e-09 wk1 = 8.781247586e-07 pk1 = -8.036475234e-13   k2 = 4.452504818e-02 lk2 = -1.613377947e-09 wk2 = -2.632996099e-07 pk2 = 1.612349128e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 6.263746314e-01 ldsub = -1.039300731e-07 wdsub = -6.633230560e-06 pdsub = 1.038637989e-11   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.699701984e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.990376632e-09 wvoff = 2.418595101e-07 pvoff = -3.987832048e-13   nfactor = {1.492059352e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.436116644e-08 wnfactor = 4.534731272e-06 pnfactor = -4.433287821e-12   eta0 = 1.030653997e-01 leta0 = -3.509075451e-08 weta0 = -2.305069136e-06 peta0 = 3.506837783e-12   etab = -7.522260139e-02 letab = 8.001307021e-11 wetab = 5.219271041e-07 petab = -7.996204747e-15   u0 = 9.698019529e-03 lu0 = -1.469720240e-10 wu0 = -1.981510912e-08 pu0 = 1.468783029e-14   ua = 1.316120392e-11 lua = 2.078860224e-17 wua = -2.106271408e-15 pua = -2.077534576e-21   ub = 3.208121026e-20 lub = -5.619352006e-26 wub = -9.426945048e-25 pub = 5.615768658e-30   uc = -6.955109697e-11 luc = -1.412099948e-18 wuc = -8.659075066e-17 puc = 1.411199480e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.333259606e+05 lvsat = -5.083180582e-03 wvsat = -7.603678806e-01 pvsat = 5.079939140e-7   a0 = 1.859769241e+00 la0 = 1.652845994e-08 wa0 = 8.462358917e-07 pa0 = -1.651792007e-12   ags = 5.247565009e-01 lags = -3.765365796e-08 wags = -5.616067375e-07 pags = 3.762964697e-12   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -5.397700691e-02 lketa = -2.522160957e-09 wketa = -1.402899920e-07 pketa = 2.520552626e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.434070907e-01 lpclm = -1.807107033e-08 wpclm = -1.058783478e-06 ppclm = 1.805954677e-12   pdiblc1 = 3.864485001e-01 lpdiblc1 = 7.272672798e-09 wpdiblc1 = 3.549235223e-07 ppdiblc1 = -7.268035160e-13   pdiblc2 = 5.100792454e-04 lpdiblc2 = -2.978654086e-11 wpdiblc2 = -3.199287121e-09 ppdiblc2 = 2.976754658e-15   pdiblcb = -6.981508827e-04 lpdiblcb = -3.193188810e-11 wpdiblcb = -7.287957379e-09 ppdiblcb = 3.191152578e-15   drout = 5.826162123e-01 ldrout = -4.631291406e-08 wdrout = -2.260179035e-06 pdrout = 4.628338124e-12   pscbe1 = 800000000.0   pscbe2 = 9.005069375e-09 lpscbe2 = -6.908664537e-17 wpscbe2 = -5.444353553e-15 ppscbe2 = 6.904259019e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.287867324e+00 lbeta0 = -2.432373010e-07 wbeta0 = 2.853976483e-06 pbeta0 = 2.430821935e-11   agidl = 1.479139429e-10 lagidl = 8.446211696e-19 wagidl = -2.573740590e-16 pagidl = -8.440825716e-23   bgidl = 1.009888412e+09 lbgidl = -2.024924373e+01 wbgidl = -9.882106772e+02 pbgidl = 2.023633119e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.572272696e-01 lkt1 = 6.434319852e-09 wkt1 = 4.764229565e-07 pkt1 = -6.430216815e-13   kt2 = -4.036919528e-02 lkt2 = 5.588370465e-10 wkt2 = 2.318049011e-09 pkt2 = -5.584806873e-14   at = 2.796473572e+05 lat = -8.883543935e-03 wat = -1.712642901e+00 pat = 8.877879077e-7   ute = -4.052831784e-01 lute = 1.990750151e-07 wute = 1.069649255e-05 pute = -1.989480689e-11   ua1 = 2.268083465e-09 lua1 = 3.968862813e-16 wua1 = 1.502206816e-14 pua1 = -3.966331949e-20   ub1 = -8.830617707e-19 lub1 = -2.241681173e-25 wub1 = -8.470418064e-24 pub1 = 2.240251697e-29   uc1 = 1.581578248e-10 luc1 = -1.153393208e-17 wuc1 = -2.122428189e-15 puc1 = 1.152657712e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.096732828e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.391677667e-09 wvth0 = -6.704539814e-08 pvth0 = 5.305320094e-14   k1 = 3.547101031e-01 lk1 = 7.739562851e-08 wk1 = 3.589975205e-07 pk1 = -2.597189815e-13   k2 = 7.197427342e-02 lk2 = -3.037398992e-08 wk2 = -2.954305201e-07 pk2 = 1.949008773e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 7.737684973e-01 ldsub = -2.583656810e-07 wdsub = 1.569194188e-06 pdsub = 1.792084304e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.731013791e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.271149516e-09 wvoff = -1.373630483e-07 pvoff = -1.443288683e-15   nfactor = {1.203943963e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.462412680e-07 wnfactor = -1.482070232e-06 pnfactor = 1.870966375e-12   eta0 = 1.463675910e-01 leta0 = -8.046170802e-08 weta0 = 2.071541574e-06 peta0 = -1.078865503e-12   etab = -1.569657760e-01 letab = 8.572846783e-08 wetab = 1.081814806e-06 petab = -5.946325419e-13   u0 = 1.138398568e-02 lu0 = -1.913485213e-09 wu0 = -2.598400744e-09 pu0 = -3.351406330e-15   ua = 4.784435631e-10 lua = -4.667226216e-16 wua = -2.763419366e-15 pua = -1.388991374e-21   ub = -2.756556127e-19 lub = 2.662454296e-25 wub = 3.375887087e-24 pub = 1.090866831e-30   uc = -6.409679862e-11 luc = -7.126977397e-18 wuc = -3.720163966e-16 puc = 4.401818042e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.083644240e+05 lvsat = -8.370660660e-02 wvsat = -7.343145546e-01 pvsat = 4.806958903e-7   a0 = 1.813205521e+00 la0 = 6.531676230e-08 wa0 = 4.917834649e-06 pa0 = -5.917911395e-12   ags = 2.880620859e-01 lags = 2.103488327e-07 wags = 4.349897085e-06 pags = -1.383186220e-12   a1 = 0.0   a2 = 8.163410947e-01 la2 = -1.712179046e-08 wa2 = -1.633067427e-06 pa2 = 1.711087224e-12   b0 = 0.0   b1 = 0.0   keta = -5.275464468e-02 lketa = -3.802921546e-09 wketa = -9.759523059e-09 pketa = 1.152887005e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.677530569e-01 lpclm = -4.358016503e-08 wpclm = -8.937474429e-07 ppclm = 1.633034045e-12   pdiblc1 = 3.697948868e-01 lpdiblc1 = 2.472191242e-08 wpdiblc1 = 2.019222879e-06 ppdiblc1 = -2.470614775e-12   pdiblc2 = 7.856911068e-04 lpdiblc2 = -3.185657589e-10 wpdiblc2 = -5.101321930e-09 ppdiblc2 = 4.969659179e-15   pdiblcb = -1.756886807e-03 lpdiblcb = 1.077385145e-09 wpdiblcb = 1.826801734e-07 ppdiblcb = -1.958527057e-13   drout = 5.468984786e-01 ldrout = -8.888765660e-09 wdrout = 1.309316683e-06 pdrout = 8.883097472e-13   pscbe1 = 7.966470932e+08 lpscbe1 = 3.513091927e+00 wpscbe1 = 3.350768723e+02 ppscbe1 = -3.510851699e-4   pscbe2 = 9.269066620e-09 lpscbe2 = -3.456963588e-16 wpscbe2 = -1.380477388e-15 ppscbe2 = 2.646231171e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 2.751125136e+00 lbeta0 = 2.414697745e-06 wbeta0 = 4.007817899e-05 pbeta0 = -1.469436943e-11   agidl = 1.958817058e-10 lagidl = -4.941480165e-17 wagidl = -6.650577560e-16 pagidl = 3.427525285e-22   bgidl = 9.940412584e+08 lbgidl = -3.644991955e+00 wbgidl = 5.954941810e+02 pbgidl = 3.642667616e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.783320628e-01 lkt1 = 2.854739459e-08 wkt1 = 1.998752925e-07 pkt1 = -3.532619528e-13   kt2 = -3.470786295e-02 lkt2 = -5.372965441e-09 wkt2 = -1.968979274e-07 pkt2 = 1.528854509e-13   at = 4.645034199e+05 lat = -2.025711051e-01 wat = -1.397716573e+00 pat = 5.578159750e-7   ute = -2.639824389e-01 lute = 5.102363275e-08 wute = -1.783686618e-05 pute = 1.000173304e-11   ua1 = 3.595855707e-09 lua1 = -9.943202802e-16 wua1 = -5.381875368e-14 pua1 = 3.246637261e-20   ub1 = -1.719809681e-18 lub1 = 6.525554249e-25 wub1 = 3.887639902e-23 pub1 = -2.720629430e-29   uc1 = 3.775330426e-10 luc1 = -2.413898009e-16 wuc1 = -1.137837795e-15 puc1 = 1.210285128e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.081333394e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.374725284e-11 wvth0 = 2.182551662e-08 pvth0 = 4.371935609e-15   k1 = 5.197901185e-01 lk1 = -1.303107693e-08 wk1 = -2.492530403e-06 pk1 = 1.302276727e-12   k2 = 6.994732204e-03 lk2 = 5.220178269e-09 wk2 = 1.012744960e-06 pk2 = -5.216849465e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.739896710e-01 ldsub = 1.540066561e-08 wdsub = 7.650466235e-06 pdsub = -1.539084492e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.629593062e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.715575527e-09 wvoff = 1.729922349e-07 pvoff = -1.714481539e-13   nfactor = {1.816790683e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.053915603e-08 wnfactor = 3.856271089e-06 pnfactor = -1.053243542e-12   eta0 = 4.174885777e-02 leta0 = -2.315418140e-08 weta0 = -4.122255420e-06 peta0 = 2.313941645e-12   etab = -4.293949384e-04 letab = -1.824829790e-11 wetab = -7.056003813e-09 petab = 1.823666133e-15   u0 = 7.717235778e-03 lu0 = 9.506871719e-11 wu0 = 8.627746939e-09 pu0 = -9.500809377e-15   ua = -4.357215007e-10 lua = 3.403414615e-17 wua = 9.100833528e-16 pua = -3.401244326e-21   ub = 2.723834647e-19 lub = -3.395667605e-26 wub = -8.277283111e-25 pub = 3.393502255e-30   uc = -7.578311593e-11 luc = -7.255049365e-19 wuc = 2.992036746e-16 puc = 7.250422965e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.572797021e+04 lvsat = -9.617310418e-05 wvsat = 1.256821825e-01 pvsat = 9.611177652e-9   a0 = 1.905621627e+00 la0 = 1.469352947e-08 wa0 = -3.205017662e-06 pa0 = -1.468415970e-12   ags = 7.938665548e-01 lags = -6.671821024e-08 wags = -1.034729201e-05 pags = 6.667566537e-12   a1 = 0.0   a2 = 7.673178107e-01 la2 = 9.731938926e-09 wa2 = 3.266134855e-06 pa2 = -9.725733064e-13   b0 = 0.0   b1 = 0.0   keta = -6.473750872e-02 lketa = 2.760991804e-09 wketa = 7.044238879e-07 pketa = -2.759231174e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.733611288e-01 lpclm = 8.125373378e-09 wpclm = 3.569861236e-06 ppclm = -8.120191990e-13   pdiblc1 = 4.432670591e-01 lpdiblc1 = -1.552430674e-08 wpdiblc1 = -5.323309172e-06 ppdiblc1 = 1.551440720e-12   pdiblc2 = 8.876357917e-04 lpdiblc2 = -3.744085086e-10 wpdiblc2 = -6.433607416e-08 ppdiblc2 = 3.741697558e-14   pdiblcb = 2.099520320e-04 wpdiblcb = -1.748620760e-7   drout = 4.959293182e-01 ldrout = 1.903086618e-08 wdrout = 6.402982523e-06 pdrout = -1.901873058e-12   pscbe1 = 8.067058136e+08 lpscbe1 = -1.996823648e+00 wpscbe1 = -6.701537446e+02 ppscbe1 = 1.995550313e-4   pscbe2 = 7.915256751e-09 lpscbe2 = 3.958868424e-16 wpscbe2 = 7.567610697e-14 ppscbe2 = -3.956343933e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.493026130e-09 lalpha0 = -7.630648883e-16 walpha0 = -1.392137825e-13 palpha0 = 7.625782971e-20   alpha1 = 9.111640222e-11 lalpha1 = 4.866212774e-18 walpha1 = 8.877932887e-16 palpha1 = -4.863109687e-22   beta0 = 7.832608366e+00 lbeta0 = -3.688117309e-07 wbeta0 = -5.403349849e-05 pbeta0 = 3.685765470e-11   agidl = 1.056716713e-10 wagidl = -3.934002799e-17   bgidl = 9.938881780e+08 lbgidl = -3.561138304e+00 wbgidl = 6.107924658e+02 pbgidl = 3.558867437e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.267952123e-01 lkt1 = 3.167962910e-10 wkt1 = -3.872316860e-07 pkt1 = -3.165942764e-14   kt2 = -4.502351865e-02 lkt2 = 2.776928650e-10 wkt2 = 1.328670847e-07 pkt2 = -2.775157859e-14   at = 9.516595301e+04 lat = -2.572741389e-04 wat = -4.263232697e-01 pat = 2.571100803e-8   ute = -1.655052166e-01 lute = -2.919727664e-09 wute = -1.107076964e-07 pute = 2.917865812e-13   ua1 = 1.659533376e-09 lua1 = 6.634868464e-17 wua1 = 1.755546046e-14 pua1 = -6.630637541e-21   ub1 = -4.093713060e-19 lub1 = -6.526995621e-26 wub1 = -2.269838586e-23 pub1 = 6.522833487e-30   uc1 = -5.237426432e-11 luc1 = -5.897325839e-18 wuc1 = -1.992801988e-15 puc1 = 5.893565233e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.078416503e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.123245834e-10 wvth0 = -2.696776170e-07 pvth0 = 9.117428123e-14   k1 = 5.335248558e-01 lk1 = -1.712093833e-08 wk1 = -3.865128296e-06 pk1 = 1.711002065e-12   k2 = 1.791124258e-03 lk2 = 6.769682625e-09 wk2 = 1.532773931e-06 pk2 = -6.765365733e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.969444487e-01 ldsub = 8.565306682e-09 wdsub = 5.356452245e-06 pdsub = -8.559844757e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.619243661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.407396233e-09 wvoff = 6.956421880e-08 pvoff = -1.406498764e-13   nfactor = {1.816691497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.056869109e-08 wnfactor = 3.866183346e-06 pnfactor = -1.056195165e-12   eta0 = -3.600844692e-02 weta0 = 3.648516622e-6   etab = -4.906771148e-04 letab = 2.167994408e-18 wetab = -9.316940175e-10 petab = -2.166611959e-22   u0 = 7.839902024e-03 lu0 = 5.854177593e-11 wu0 = -3.631055432e-09 pu0 = -5.850444501e-15   ua = -4.156218658e-10 lua = 2.804897739e-17 wua = -1.098598418e-15 pua = -2.803109112e-21   ub = 2.501698715e-19 lub = -2.734202331e-26 wub = 1.392214501e-24 pub = 2.732458785e-30   uc = -8.087943093e-11 luc = 7.920502627e-19 wuc = 8.085101928e-16 puc = -7.915451880e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.757705730e+04 lvsat = -6.467850102e-04 wvsat = -5.910861316e-02 pvsat = 6.463725683e-8   a0 = 1.912010217e+00 la0 = 1.279116724e-08 wa0 = -3.843469222e-06 pa0 = -1.278301057e-12   ags = 3.134834868e-01 lags = 7.632785785e-08 wags = 3.766038172e-05 pags = -7.627918510e-12   a1 = 0.0   a2 = 7.816984453e-01 la2 = 5.449745456e-09 wa2 = 1.828988418e-06 pa2 = -5.446270262e-13   b0 = 0.0   b1 = 0.0   keta = -5.563944227e-02 lketa = 5.181506729e-11 wketa = -2.048025913e-07 pketa = -5.178202586e-15   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.960454667e-01 lpclm = 1.370544663e-09 wpclm = 1.302873982e-06 ppclm = -1.369670694e-13   pdiblc1 = 3.990851626e-01 lpdiblc1 = -2.368042522e-09 wpdiblc1 = -9.079369183e-07 ppdiblc1 = 2.366532468e-13   pdiblc2 = -2.081112101e-04 lpdiblc2 = -4.812244520e-11 wpdiblc2 = 4.516875242e-08 ppdiblc2 = 4.809175848e-15   pdiblcb = -3.628799332e-02 lpdiblcb = 1.086817568e-08 wpdiblcb = 3.472605058e-06 ppdiblcb = -1.086124526e-12   drout = 5.654052296e-01 ldrout = -1.657323355e-09 wdrout = -5.401782841e-07 pdrout = 1.656266513e-13   pscbe1 = 7.999751827e+08 lpscbe1 = 7.389970407e-03 wpscbe1 = 2.480147081e+00 ppscbe1 = -7.385257970e-7   pscbe2 = 1.125473216e-08 lpscbe2 = -5.985254465e-16 wpscbe2 = -2.580584819e-13 ppscbe2 = 5.981437788e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.377503366e-09 lalpha0 = 9.170703233e-17 walpha0 = 1.476561192e-13 palpha0 = -9.164855258e-21   alpha1 = 1.074583140e-10 walpha1 = -7.453557961e-16   beta0 = 6.481398941e+00 lbeta0 = 3.354465542e-08 wbeta0 = 8.100128000e-05 pbeta0 = -3.352326466e-12   agidl = 1.056716713e-10 wagidl = -3.934002799e-17   bgidl = 1.019536931e+09 lbgidl = -1.119869583e+01 wbgidl = -1.952447297e+03 pbgidl = 1.119155464e-3   cgidl = 2.390949645e+02 lcgidl = 1.813599694e-05 wcgidl = 6.086619756e-03 pcgidl = -1.812443198e-9   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.307799964e-01 lkt1 = 1.503365398e-09 wkt1 = 1.099262941e-08 pkt1 = -1.502406732e-13   kt2 = -4.766196413e-02 lkt2 = 1.063355965e-09 wkt2 = 3.965433835e-07 pkt2 = -1.062677885e-13   at = 9.132686249e+04 lat = 8.859110399e-04 wat = -4.265902913e-02 pat = -8.853461121e-8   ute = -2.036903229e-01 lute = 8.450842356e-09 wute = 3.705367943e-06 pute = -8.445453423e-13   ua1 = 1.682025175e-09 lua1 = 5.965118928e-17 wua1 = 1.530771485e-14 pua1 = -5.961315091e-21   ub1 = -4.311756146e-19 lub1 = -5.877717822e-26 wub1 = -2.051934541e-23 pub1 = 5.873969718e-30   uc1 = -5.645680963e-11 luc1 = -4.681645908e-18 wuc1 = -1.584807792e-15 puc1 = 4.678660516e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.088591948e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.510278560e-09 wvth0 = 7.472180113e-07 pvth0 = -1.509315486e-13   k1 = 5.107715443e-01 lk1 = -1.282931870e-08 wk1 = -1.591248079e-06 pk1 = 1.282113770e-12   k2 = -3.022497284e-04 lk2 = 7.787343887e-09 wk2 = 1.741977840e-06 pk2 = -7.782378054e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.979910879e-01 ldsub = 3.342588772e-08 wdsub = 1.524547827e-05 pdsub = -3.340457270e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.624546845e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.642246018e-09 wvoff = 1.225622422e-07 pvoff = -1.641198791e-13   nfactor = {2.169286295e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.494890585e-08 wnfactor = -3.137081224e-05 pnfactor = 7.490111243e-12   eta0 = -1.801757916e-01 leta0 = 3.528856178e-08 weta0 = 1.805605782e-05 peta0 = -3.526605897e-12   etab = -1.930138233e-02 letab = 4.604390370e-09 wetab = 1.878939306e-06 petab = -4.601454243e-13   u0 = 8.841579544e-03 lu0 = -1.822745705e-10 wu0 = -1.037349325e-07 pu0 = 1.821583376e-14   ua = -7.905413624e-11 lua = -5.224095160e-17 wua = -3.473390912e-14 pua = 5.220763859e-21   ub = -3.117057615e-20 lub = 3.948241130e-26 wub = 2.950831874e-23 pub = -3.945723416e-30   uc = -7.957484394e-11 luc = 5.318346988e-19 wuc = 6.781346849e-16 puc = -5.314955584e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.734342161e+04 lvsat = 4.257630328e-03 wvsat = 1.962964697e+00 pvsat = -4.254915322e-7   a0 = 1.961791845e+00 la0 = 1.560538621e-09 wa0 = -8.818457594e-06 pa0 = -1.559543497e-13   ags = 6.485854859e-01 wags = 4.171550598e-6   a1 = 0.0   a2 = 8.372605790e-01 la2 = -7.743733760e-09 wa2 = -3.723681866e-06 pa2 = 7.738795736e-13   b0 = 1.125199427e-24 lb0 = -2.754206898e-31 wb0 = -1.124481910e-28 pb0 = 2.752450595e-35   b1 = 0.0   keta = -1.989339662e-02 lketa = -8.694056036e-09 wketa = -3.777127702e-06 pketa = 8.688512010e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.618317068e-01 lpclm = 9.847508422e-09 wpclm = 4.722068229e-06 ppclm = -9.841228863e-13   pdiblc1 = 2.664210246e-01 lpdiblc1 = 2.992808286e-08 wpdiblc1 = 1.235001715e-05 ppdiblc1 = -2.990899832e-12   pdiblc2 = -3.238752328e-03 lpdiblc2 = 6.901111129e-10 wpdiblc2 = 3.480396062e-07 ppdiblc2 = -6.896710429e-14   pdiblcb = 1.497212350e-02 lpdiblcb = -8.678725116e-10 wpdiblcb = -1.650137869e-06 ppdiblcb = 8.673190867e-14   drout = 7.796742867e-01 ldrout = -5.422872623e-08 wdrout = -2.195342048e-05 pdrout = 5.419414565e-12   pscbe1 = 8.000622289e+08 lpscbe1 = -1.336521603e-02 wpscbe1 = -6.218923663e+00 ppscbe1 = 1.335669330e-6   pscbe2 = 8.751261867e-09 lpscbe2 = -3.040948681e-17 wpscbe2 = -7.871094210e-15 ppscbe2 = 3.039009529e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -5.715221550e-09 lalpha0 = 1.160316560e-15 walpha0 = 5.811513300e-13 palpha0 = -1.159576650e-19   alpha1 = 1.074583140e-10 walpha1 = -7.453557961e-16   beta0 = 5.380643155e+00 lbeta0 = 3.054857602e-07 wbeta0 = 1.910066656e-04 pbeta0 = -3.052909581e-11   agidl = 1.056716713e-10 wagidl = -3.934002799e-17   bgidl = 9.100084584e+08 lbgidl = 1.477532082e+01 wbgidl = 8.993415575e+03 pbgidl = -1.476589889e-3   cgidl = 4.527182679e+02 lcgidl = -3.280006599e-05 wcgidl = -1.526208825e-02 pcgidl = 3.277915004e-9   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.299731666e-01 lkt1 = 1.418077390e-09 wkt1 = -6.963890259e-08 pkt1 = -1.417173110e-13   kt2 = -3.631482942e-02 lkt2 = -1.634775299e-09 wkt2 = -7.374465027e-07 pkt2 = 1.633732836e-13   at = 9.081810355e+04 lat = 1.076562531e-03 wat = 8.184422798e-03 pat = -1.075876029e-7   ute = -2.269573520e-01 lute = 1.477675850e-08 wute = 6.030587161e-06 pute = -1.476733566e-12   ua1 = 1.962749505e-09 lua1 = -4.611038739e-18 wua1 = -1.274681693e-14 pua1 = 4.608098372e-22   ub1 = -7.490634351e-19 lub1 = 1.464697501e-26 wub1 = 1.124916556e-23 pub1 = -1.463763493e-30   uc1 = -9.155673900e-11 luc1 = 3.560524395e-18 wuc1 = 1.922946892e-15 puc1 = -3.558253920e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.094013643e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.108886765e-07 wvth0 = -7.687823004e-09 pvth0 = 7.691495862e-13   k1 = 4.350917301e-01 lk1 = 1.480796990e-07 wk1 = 1.026624677e-08 pk1 = -1.027115147e-12   k2 = 3.861023817e-02 lk2 = 2.159309455e-08 wk2 = 1.497031927e-09 pk2 = -1.497747134e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.742543315e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.932284296e-07 wvoff = 4.112805124e-08 pvoff = -4.114770017e-12   nfactor = {1.469021010e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.298786098e-05 wnfactor = 9.004379854e-07 pnfactor = -9.008681696e-11   eta0 = 0.08   etab = -0.07   u0 = 9.215150546e-03 lu0 = 1.325107308e-08 wu0 = 9.186862688e-10 pu0 = -9.191251712e-14   ua = -8.495126258e-11 lua = 3.238975939e-15 wua = 2.245556041e-16 pua = -2.246628856e-20   ub = 9.992607462e-20 lub = -2.322543527e-24 wub = -1.610200800e-25 pub = 1.610970073e-29   uc = -7.883729334e-11 luc = 1.167154680e-16 wuc = 8.091789789e-18 puc = -8.095655641e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.754531650e+05 lvsat = 2.455856221e+00 wvsat = 1.702625421e-01 pvsat = -1.703438850e-5   a0 = 1.679650653e+00 la0 = -8.170366789e-06 wa0 = -5.664449767e-07 pa0 = 5.667155958e-11   ags = 3.609097476e-01 lags = -9.532146567e-06 wags = -6.608560764e-07 pags = 6.611718004e-11   a1 = 0.0   a2 = 8.762955994e-01 la2 = 1.237534956e-05 wa2 = 8.579730595e-07 pa2 = -8.583829561e-11   b0 = 0.0   b1 = 0.0   keta = -3.600581574e-02 lketa = 2.284764399e-06 wketa = 1.584008833e-07 pketa = -1.584765593e-11   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.373215098e-01 lpclm = -6.186138797e-06 wpclm = -4.288800414e-07 ppclm = 4.290849388e-11   pdiblc1 = 0.39   pdiblc2 = 1.486829619e-03 lpdiblc2 = 2.141792534e-07 wpdiblc2 = 1.484887586e-08 ppdiblc2 = -1.485596991e-12   pdiblcb = -1.932410293e-03 lpdiblcb = 1.837543721e-07 wpdiblcb = 1.273954324e-08 ppdiblcb = -1.274562956e-12   drout = 0.56   pscbe1 = 7.293227697e+08 lpscbe1 = 1.716055485e+03 wpscbe1 = 1.189727505e+02 ppscbe1 = -1.190295897e-2   pscbe2 = 9.566796900e-09 lpscbe2 = -6.183392694e-15 wpscbe2 = -4.286896562e-16 ppscbe2 = 4.288944627e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 3.316586945e-10 lalpha0 = -2.317693695e-14 walpha0 = -1.606838450e-15 palpha0 = 1.607606117e-19   alpha1 = 3.831996208e-11 lalpha1 = 6.170950555e-15 walpha1 = 4.278270528e-16 palpha1 = -4.280314471e-20   beta0 = 3.816634675e+00 lbeta0 = 9.762205917e-05 wbeta0 = 6.768059067e-06 pbeta0 = -6.771292508e-10   agidl = 1.0e-10   bgidl = 1.337499634e+09 lbgidl = -1.831424881e+04 wbgidl = -1.269712181e+03 pbgidl = 1.270318786e-1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.355049707e-01 lkt1 = -6.187984178e-07 wkt1 = -4.290079801e-08 pkt1 = 4.292129387e-12   kt2 = -0.037961   at = 0.0   ute = -3.316284416e-01 lute = 3.098323678e-06 wute = 2.148042957e-07 pute = -2.149069184e-11   ua1 = 2.2116e-9   ub1 = -8.721213168e-19 lub1 = 7.856883511e-24 wub1 = 5.447114324e-25 pub1 = -5.449716683e-29   uc1 = 1.1985e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.099544864e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.067800992e-8   k1 = 4.424780710e-01 wk1 = -4.096712684e-8   k2 = 3.968732001e-02 wk2 = -5.973857655e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.446635949e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = -1.641201629e-7   nfactor = {2.116866518e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -3.593168760e-6   eta0 = 0.08   etab = -0.07   u0 = 9.876125296e-03 wu0 = -3.665987947e-9   ua = 7.661160111e-11 wua = -8.960819009e-16   ub = -1.592436400e-20 wub = 6.425454396e-25   uc = -7.301542692e-11 wuc = -3.229002635e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.979533538e+05 wvsat = -6.794271868e-1   a0 = 1.272105836e+00 wa0 = 2.260380423e-6   ags = -1.145617981e-01 wags = 2.637124874e-6   a1 = 0.0   a2 = 1.493588519e+00 wa2 = -3.423713842e-6   b0 = 0.0   b1 = 0.0   keta = 7.796016795e-02 wketa = -6.320936196e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.712483338e-01 wpclm = 1.711431982e-6   pdiblc1 = 0.39   pdiblc2 = 1.217027222e-02 wpdiblc2 = -5.925396055e-8   pdiblcb = 7.233413451e-03 wpdiblcb = -5.083673672e-8   drout = 0.56   pscbe1 = 8.149210710e+08 wpscbe1 = -4.747569262e+2   pscbe2 = 9.258364034e-09 wpscbe2 = 1.710672257e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -8.244265541e-10 walpha0 = 6.412037046e-15   alpha1 = 3.461322034e-10 walpha1 = -1.707230065e-15   beta0 = 8.686105685e+00 wbeta0 = -2.700772157e-5   agidl = 1.0e-10   bgidl = 4.239693885e+08 wbgidl = 5.066745537e+3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.663711600e-01 wkt1 = 1.711942518e-7   kt2 = -0.037961   at = 0.0   ute = -1.770814319e-01 wute = -8.571696187e-7   ua1 = 2.2116e-9   ub1 = -4.802133115e-19 wub1 = -2.173653415e-24   uc1 = 1.1985e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.104158953e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.713315161e-08 wvth0 = 1.892547934e-08 pvth0 = 9.458172179e-14   k1 = 6.139589363e-01 lk1 = -1.380039421e-06 wk1 = -1.182084835e-06 pk1 = 9.183458565e-12   k2 = -2.799883308e-02 lk2 = 5.447229307e-07 wk2 = 4.420044048e-07 pk2 = -3.605228261e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.563423265e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.398780408e-08 wvoff = -8.855229213e-08 pvoff = -6.081532214e-13   nfactor = {1.575456415e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.357146697e-06 wnfactor = 5.931626695e-07 pnfactor = -3.369065342e-11   eta0 = 0.08   etab = -0.07   u0 = 7.543599058e-03 lu0 = 1.877164635e-08 wu0 = 1.144504480e-08 pu0 = -1.216101915e-13   ua = -5.679814196e-10 lua = 5.187539597e-15 wua = 3.261478696e-15 pua = -3.345911223e-20   ub = 4.458446464e-19 lub = -3.716213097e-24 wub = -2.180915838e-24 pub = 2.272258109e-29   uc = -1.288331838e-10 luc = 4.492087486e-16 wuc = 3.039645469e-16 puc = -2.706101148e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.965941337e+05 lvsat = -7.938388030e-01 wvsat = -8.422274709e-01 pvsat = 1.310180056e-6   a0 = 6.183607608e-01 la0 = 5.261193271e-06 wa0 = 4.897995456e-06 pa0 = -2.122693232e-11   ags = -6.442177027e-01 lags = 4.262551548e-06 wags = 4.531583777e-06 pags = -1.524617900e-11   a1 = 0.0   a2 = 2.195461086e+00 la2 = -5.648512496e-06 wa2 = -6.888319665e-06 pa2 = 2.788236813e-11   b0 = 0.0   b1 = 0.0   keta = 2.223657241e-01 lketa = -1.162143425e-06 wketa = -1.337436762e-06 pketa = 5.676442910e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -9.849126693e-01 lpclm = 6.548187497e-06 wpclm = 3.443304881e-06 ppclm = -1.393772341e-11   pdiblc1 = 0.39   pdiblc2 = 2.334509515e-02 lpdiblc2 = -8.993246063e-08 wpdiblc2 = -1.146583084e-07 ppdiblc2 = 4.458817258e-13   pdiblcb = 9.639393160e-03 lpdiblcb = -1.936278335e-08 wpdiblcb = -6.278495665e-08 ppdiblcb = 9.615658568e-14   drout = 0.56   pscbe1 = 6.401950268e+08 lpscbe1 = 1.406155890e+03 wpscbe1 = 3.614882892e+02 ppscbe1 = -6.729913339e-3   pscbe2 = 9.825805884e-09 lpscbe2 = -4.566644332e-15 wpscbe2 = 1.666149846e-15 ppscbe2 = 3.583063458e-22   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.759894228e-09 lalpha0 = 7.528433358e-15 walpha0 = 1.290065786e-14 palpha0 = -5.221896037e-20   alpha1 = 5.952041482e-10 lalpha1 = -2.004474971e-15 walpha1 = -3.434850859e-15 palpha1 = 1.390350344e-20   beta0 = 1.372465216e+01 lbeta0 = -4.054908838e-05 wbeta0 = -6.563449912e-05 pbeta0 = 3.108596147e-10   agidl = 9.292715563e-09 lagidl = -7.398090649e-14 wagidl = -6.408104268e-14 pagidl = 5.157098133e-19   bgidl = 2.406156110e+09 lbgidl = -1.595219274e+04 wbgidl = -7.598102948e+03 pbgidl = 1.019238510e-1   cgidl = 300.0   egidl = 6.239518307e-01 legidl = -4.216646444e-06 wegidl = -3.634251454e-06 pegidl = 2.924763800e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.384389309e-01 lkt1 = -2.247922950e-07 wkt1 = 5.304528575e-08 pkt1 = 9.508362952e-13   kt2 = -4.604989928e-02 lkt2 = 6.509764143e-08 wkt2 = 7.284697979e-08 pkt2 = -5.862561028e-13   at = -4.640542657e+05 lat = 3.734604318e+00 wat = 1.376210244e+00 pat = -1.107543039e-5   ute = -2.286690795e+00 lute = 1.697766149e-05 wute = 1.375865438e-05 pute = -1.176248630e-10   ua1 = -4.881515119e-09 lua1 = 5.708379453e-14 wua1 = 4.774794702e-14 pua1 = -3.842647344e-19   ub1 = 4.287650512e-18 lub1 = -3.837069528e-23 wub1 = -3.402172932e-23 pub1 = 2.563061491e-28   uc1 = -8.794039289e-11 luc1 = 1.672250329e-15 wuc1 = 1.321466735e-15 puc1 = -1.063486695e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.133317561e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.551606369e-07 wvth0 = 2.529705108e-07 pvth0 = -8.527799054e-13   k1 = 1.434459846e-01 lk1 = 5.244911420e-07 wk1 = 1.522682782e-06 pk1 = -1.764832175e-12   k2 = 1.477164608e-01 lk2 = -1.665330429e-07 wk2 = -5.581784614e-07 pk2 = 4.432869401e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.303773026e+00 ldsub = -3.010625861e-06 wdsub = -3.671436212e-06 pdsub = 1.486114771e-11   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.642719863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.260852829e-07 wvoff = -6.763426337e-08 pvoff = -6.928246952e-13   nfactor = {1.895827954e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.060354790e-06 wnfactor = -4.743894398e-06 pnfactor = -1.208744725e-11   eta0 = 3.623013694e-01 leta0 = -1.142692425e-06 weta0 = -1.393505053e-06 peta0 = 5.640594916e-12   etab = -3.167917632e-01 letab = 9.989575291e-07 wetab = 1.218221399e-06 petab = -4.931086122e-12   u0 = 1.498354271e-02 lu0 = -1.134357155e-08 wu0 = -2.599082191e-08 pu0 = 2.992177383e-14   ua = 9.087341851e-10 lua = -7.898729094e-16 wua = -3.384517279e-15 pua = -6.557615876e-21   ub = -2.117680564e-19 lub = -1.054344839e-24 wub = -8.881181806e-26 pub = 1.425421473e-29   uc = 7.082025245e-11 luc = -3.589434395e-16 wuc = -9.628152048e-16 puc = 2.421538261e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.934158880e+05 lvsat = -3.761964794e-01 wvsat = -6.750673245e-01 pvsat = 6.335533948e-7   a0 = 1.606562303e+00 la0 = 1.261175772e-06 wa0 = 1.777296794e-06 pa0 = -8.595046297e-12   ags = 3.629524229e-01 lags = 1.857534926e-07 wags = -1.324518736e-07 pags = 3.632787907e-12   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.720740318e-02 lketa = 9.093894062e-08 wketa = 2.371477321e-07 pketa = -6.971208419e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.714890908e-01 lpclm = 1.462555863e-06 wpclm = 2.674751443e-06 ppclm = -1.082679202e-11   pdiblc1 = 0.39   pdiblc2 = 1.958983320e-03 lpdiblc2 = -3.366291825e-09 wpdiblc2 = -8.608706273e-09 ppdiblc2 = 1.661679743e-14   pdiblcb = 1.139832103e-02 lpdiblcb = -2.648252763e-08 wpdiblcb = -7.895046738e-08 ppdiblcb = 1.615909359e-13   drout = 0.56   pscbe1 = 1.178310626e+09 lpscbe1 = -7.720149809e+02 wpscbe1 = -2.624050273e+03 ppscbe1 = 5.354875015e-3   pscbe2 = 9.711142554e-09 lpscbe2 = -4.102512971e-15 wpscbe2 = -3.300385212e-15 ppscbe2 = 2.046172279e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.801102460e-03 lalpha0 = -1.133823210e-08 walpha0 = -1.942909582e-08 palpha0 = 7.864460835e-14   alpha1 = -1.527073121e-10 lalpha1 = 1.022902340e-15 walpha1 = 1.752836545e-15 palpha1 = -7.095087945e-21   beta0 = 6.822857684e+01 lbeta0 = -2.611687121e-04 wbeta0 = -4.504031476e-04 pbeta0 = 1.868316531e-9   agidl = -1.830417317e-08 lagidl = 3.772508979e-14 wagidl = 1.282546004e-13 pagidl = -2.628215945e-19   bgidl = -3.285688709e+09 lbgidl = 7.087114421e+03 wbgidl = 2.972653117e+04 pbgidl = -4.915786984e-2   cgidl = 300.0   egidl = -9.479036614e-01 legidl = 2.145870920e-06 wegidl = 7.268502909e-06 pegidl = -1.488425854e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.884919984e-01 lkt1 = 3.825887605e-07 wkt1 = 7.887986367e-07 pkt1 = -2.027327725e-12   kt2 = -2.959136871e-02 lkt2 = -1.522787162e-09 wkt2 = -5.081938538e-08 pkt2 = -8.568248150e-14   at = 7.393921732e+05 lat = -1.136676091e+00 wat = -2.089004686e+00 pat = 2.950979967e-6   ute = 4.281821328e+00 lute = -9.610197668e-06 wute = -3.270331292e-05 pute = 7.044272670e-11   ua1 = 1.779649922e-08 lua1 = -3.471170498e-14 wua1 = -1.025242235e-13 pua1 = 2.240032005e-19   ub1 = -1.143012074e-17 lub1 = 2.525130624e-23 wub1 = 7.021593664e-23 pub1 = -1.656244692e-28   uc1 = 1.052975756e-09 luc1 = -2.945921535e-15 wuc1 = -4.868004757e-15 puc1 = 1.441872102e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.043507227e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.875072053e-08 wvth0 = -1.883632782e-07 pvth0 = 5.097239444e-14   k1 = 3.438755816e-01 lk1 = 1.140564239e-07 wk1 = 1.412396612e-06 pk1 = -1.538990915e-12   k2 = 1.023501676e-01 lk2 = -7.363308192e-08 wk2 = -6.643880538e-07 pk2 = 6.607802882e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -1.767772157e+00 ldsub = 3.279207576e-06 wdsub = 9.973127006e-06 pdsub = -1.307984773e-11   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.158430313e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.661069875e-07 wvoff = -7.873794849e-07 pvoff = 7.810515757e-13   nfactor = {5.413710842e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.143477841e-06 wnfactor = -2.266675329e-05 pnfactor = 2.461453511e-11   eta0 = -6.304968526e-01 leta0 = 8.903349535e-07 weta0 = 2.783088832e-06 peta0 = -2.912129626e-12   etab = -4.314104042e-01 letab = 1.233670717e-06 wetab = 2.992528340e-06 petab = -8.564467518e-12   u0 = 1.221957100e-02 lu0 = -5.683579383e-09 wu0 = -3.730517510e-08 pu0 = 5.309102342e-14   ua = 1.562850384e-09 lua = -2.129355709e-15 wua = -1.285527509e-14 pua = 1.283636520e-20   ub = -1.515888443e-18 lub = 1.616200284e-24 wub = 9.794382136e-24 pub = -5.984342765e-30   uc = -1.280980627e-10 luc = 4.839651337e-17 wuc = 3.195045866e-16 puc = -2.043641496e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.018225595e+04 lvsat = 3.998027147e-02 wvsat = -4.611131357e-01 pvsat = 1.954233558e-7   a0 = 1.182406685e+00 la0 = 2.129751043e-06 wa0 = 5.544579729e-06 pa0 = -1.630959411e-11   ags = -9.848666318e-01 lags = 2.945783657e-06 wags = 9.909489543e-06 pags = -1.693084868e-11   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 2.954023652e-02 lketa = -1.481339573e-07 wketa = -7.195849684e-07 pketa = 1.262052464e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.571468923e-01 lpclm = 5.848295836e-08 wpclm = -3.234955529e-06 ppclm = 1.274958173e-12   pdiblc1 = 5.389411732e-01 lpdiblc1 = -3.049980110e-07 wpdiblc1 = -7.028010372e-07 ppdiblc1 = 1.439178394e-12   pdiblc2 = 1.947219937e-04 lpdiblc2 = 2.465184130e-10 wpdiblc2 = -1.011896061e-09 ppdiblc2 = 1.060239395e-15   pdiblcb = -6.292190551e-02 lpdiblcb = 1.257085743e-07 wpdiblcb = 4.243104406e-07 ppdiblcb = -8.689741700e-13   drout = -1.228382711e-01 ldrout = 1.398299141e-06 wdrout = 2.633016927e-06 pdrout = -5.391826237e-12   pscbe1 = 8.026800621e+08 lpscbe1 = -2.808102096e+00 wpscbe1 = -1.858953269e+01 ppscbe1 = 1.947764762e-5   pscbe2 = 6.517198490e-09 lpscbe2 = 2.437965835e-15 wpscbe2 = 1.181209609e-14 ppscbe2 = -1.048523862e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -5.565622884e-03 lalpha0 = 5.794938887e-09 walpha0 = 3.860445224e-08 palpha0 = -4.019504054e-14   alpha1 = 3.468116000e-10 walpha1 = -1.711942518e-15   beta0 = -8.085247603e+01 lbeta0 = 4.411574095e-05 wbeta0 = 6.003433825e-04 pbeta0 = -2.833759451e-10   agidl = 1.374840824e-10 lagidl = -3.927488439e-17 wagidl = -1.850301268e-16 pagidl = 1.938699411e-22   bgidl = -1.154447506e+08 lbgidl = 5.951680990e+02 wbgidl = 6.817361219e+03 pbgidl = -2.245044346e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.531917529e-01 lkt1 = -9.925319990e-08 wkt1 = -2.451915234e-07 pkt1 = 9.005147505e-14   kt2 = -1.108277537e-02 lkt2 = -3.942422189e-08 wkt2 = -2.008193539e-07 pkt2 = 2.214837041e-13   at = 1.273251157e+05 lat = 1.166995275e-01 wat = -6.561004955e-01 pat = 1.671458901e-8   ute = 5.755912372e-01 lute = -2.020672343e-06 wute = 3.892920036e-06 pute = -4.498124237e-12   ua1 = 3.069146085e-09 lua1 = -4.553399403e-15 wua1 = 9.465711974e-15 pua1 = -5.326989513e-21   ub1 = -1.000405162e-19 lub1 = 2.049851216e-24 wub1 = -1.390163515e-23 pub1 = 6.629391309e-30   uc1 = -7.019438440e-10 luc1 = 6.477589484e-16 wuc1 = 3.843436529e-15 puc1 = -3.420350663e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.069236841e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.791874189e-09 wvth0 = -2.577639461e-07 pvth0 = 1.236886792e-13   k1 = 4.342367483e-01 lk1 = 1.937825249e-08 wk1 = -1.926177407e-07 pk1 = 1.427029986e-13   k2 = 4.486698230e-03 lk2 = 2.890581472e-08 wk2 = 1.726789585e-07 pk2 = -2.162776006e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.758410209e+00 ldsub = -4.154381524e-07 wdsub = -5.260509163e-06 pdsub = 2.881575407e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.474978341e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.059956241e-08 wvoff = 3.786680238e-07 pvoff = -4.407038527e-13   nfactor = {-2.345508273e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.986437967e-06 wnfactor = 2.313775395e-05 pnfactor = -2.337828245e-11   eta0 = 5.538851040e-01 leta0 = -3.506308510e-07 weta0 = -7.550944402e-07 peta0 = 7.950903514e-13   etab = 1.566760866e+00 letab = -8.599631857e-07 wetab = -1.087435309e-05 petab = 5.964904167e-12   u0 = 9.827439349e-03 lu0 = -3.177163647e-09 wu0 = 8.198165757e-09 pu0 = 5.413760460e-15   ua = -2.812587005e-10 lua = -1.971443127e-16 wua = 2.506051785e-15 pua = -3.258849067e-21   ub = 6.442161211e-19 lub = -6.471032749e-25 wub = -3.004556669e-24 pub = 7.426065342e-30   uc = -1.441209728e-10 luc = 6.518491800e-17 wuc = 1.830498411e-16 puc = -6.139027862e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.744794356e+05 lvsat = -1.531217060e-01 wvsat = -1.192903614e+00 pvsat = 9.621751238e-7   a0 = 6.050057499e+00 la0 = -2.970451789e-06 wa0 = -2.446995362e-05 pa0 = 1.513888357e-11   ags = 3.251405260e+00 lags = -1.492876124e-06 wags = -1.620453867e-05 pags = 1.043077723e-11   a1 = 0.0   a2 = 1.247398428e-01 la2 = 7.075207112e-07 wa2 = 3.164039307e-06 pa2 = -3.315201285e-12   b0 = 0.0   b1 = 0.0   keta = -2.046773120e-01 lketa = 9.727333460e-08 wketa = 1.044011343e-06 pketa = -5.857996618e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.504097511e-01 lpclm = 5.894294664e-07 wpclm = 6.137961495e-07 ppclm = -2.757667617e-12   pdiblc1 = 1.378932118e+00 lpdiblc1 = -1.185119524e-06 wpdiblc1 = -4.980387078e-06 ppdiblc1 = 5.921126108e-12   pdiblc2 = 2.292707366e-03 lpdiblc2 = -1.951698210e-09 wpdiblc2 = -1.555433633e-08 ppdiblc2 = 1.629744475e-14   pdiblcb = 1.469498995e-01 lpdiblcb = -9.418985618e-08 wpdiblcb = -8.487845962e-07 ppdiblcb = 4.649429822e-13   drout = 8.272671269e-01 ldrout = 4.028024572e-07 wdrout = -6.353853067e-07 pdrout = -1.967276087e-12   pscbe1 = 9.559101664e+08 lpscbe1 = -1.633587746e+02 wpscbe1 = -7.696087526e+02 ppscbe1 = 8.063768108e-4   pscbe2 = 8.950009485e-09 lpscbe2 = -1.110727058e-16 wpscbe2 = 8.325769220e-16 ppscbe2 = 1.018827082e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -7.316337109e-05 lalpha0 = 4.007712037e-11 walpha0 = 5.074788094e-10 palpha0 = -2.779842048e-16   alpha1 = 6.172060484e-10 lalpha1 = -2.833125432e-16 walpha1 = -3.587461143e-15 palpha1 = 1.965121528e-21   beta0 = -9.091879976e+01 lbeta0 = 5.466298330e-05 wbeta0 = 6.897945095e-04 pbeta0 = -3.771005996e-10   agidl = 1.0e-10   bgidl = -3.446089029e+08 lbgidl = 8.352805687e+02 wbgidl = 9.880682267e+03 pbgidl = -5.454715558e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.039606534e-01 lkt1 = -4.605881520e-08 wkt1 = -3.159820576e-07 pkt1 = 1.642240270e-13   kt2 = -7.051301275e-02 lkt2 = 2.284529508e-08 wkt2 = 5.145489847e-08 pkt2 = -4.284295071e-14   at = 4.851875060e+05 lat = -2.582597385e-01 wat = -1.541186194e+00 pat = 9.440852565e-7   ute = -2.714653968e+00 lute = 1.426764328e-06 wute = -8.384398937e-07 pute = 4.592764128e-13   ua1 = -5.640292455e-09 lua1 = 4.572132563e-15 wua1 = 1.024531276e-14 pua1 = -6.143835728e-21   ub1 = 6.604416588e-18 lub1 = -4.974911327e-24 wub1 = -1.886236560e-23 pub1 = 1.182712066e-29   uc1 = 7.472257745e-11 luc1 = -1.660127113e-16 wuc1 = 9.625258430e-16 puc1 = -4.018044682e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.047952825e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.345072581e-08 wvth0 = -2.097098547e-07 pvth0 = 9.736584928e-14   k1 = 1.777379293e-01 lk1 = 1.598818931e-07 wk1 = -1.199770628e-07 pk1 = 1.029122513e-13   k2 = 2.093729928e-01 lk2 = -8.332577530e-08 wk2 = -3.909976070e-07 pk2 = 9.249033006e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.489598722e+00 ldsub = -2.681899402e-07 wdsub = -7.812801665e-07 pdsub = 4.279657432e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.234173707e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.273531866e-08 wvoff = -8.023638478e-07 pvoff = 2.062358808e-13   nfactor = {7.593227879e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.457753228e-06 wnfactor = -3.621043743e-05 pnfactor = 9.131173080e-12   eta0 = -7.725447526e-01 leta0 = 3.759542637e-07 weta0 = 1.525873978e-06 peta0 = -4.543671238e-13   etab = -6.178572161e-03 letab = 1.653714950e-09 wetab = 3.282162321e-08 petab = -9.773458851e-15   u0 = 3.746664996e-03 lu0 = 1.537325244e-10 wu0 = 3.616854705e-08 pu0 = -9.907715154e-15   ua = 1.030703908e-09 lua = -9.158046305e-16 wua = -9.261383492e-15 pua = 3.187057792e-21   ub = -3.329073129e-18 lub = 1.529365244e-24 wub = 2.415281016e-23 pub = -7.450061274e-30   uc = -9.496408232e-11 luc = 3.825800232e-17 wuc = 4.322473076e-16 puc = -1.978944208e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.195765802e+05 lvsat = 6.273232810e-02 wvsat = 1.341635215e+00 pvsat = -4.261818829e-7   a0 = 3.321461542e-01 la0 = 1.616770981e-07 wa0 = 7.708973267e-06 pa0 = -2.487928103e-12   ags = -2.603195334e+00 lags = 1.714127716e-06 wags = 1.321551737e-05 pags = -5.684793965e-12   a1 = 0.0   a2 = 2.150520314e+00 la2 = -4.021511866e-07 wa2 = -6.328078614e-06 pa2 = 1.884343609e-12   b0 = 0.0   b1 = 0.0   keta = 6.977723432e-03 lketa = -1.866600242e-08 wketa = 2.069903998e-07 pketa = -1.273005144e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.236258247e+00 lpclm = -3.888136936e-07 wpclm = -7.964378970e-06 ppclm = 1.941242259e-12   pdiblc1 = -2.322923824e+00 lpdiblc1 = 8.426646152e-07 wpdiblc1 = 1.386363255e-05 ppdiblc1 = -4.401156743e-12   pdiblc2 = -1.269670843e-02 lpdiblc2 = 6.259129026e-09 wpdiblc2 = 2.988808891e-08 ppdiblc2 = -8.594779735e-15   pdiblcb = -0.025   drout = 2.407568336e+00 ldrout = -4.628470379e-07 wdrout = -6.856589209e-06 pdrout = 1.440543880e-12   pscbe1 = 4.881796672e+08 lpscbe1 = 9.285229961e+01 wpscbe1 = 1.539217505e+03 ppscbe1 = -4.583404926e-4   pscbe2 = 1.797497496e-08 lpscbe2 = -5.054723169e-15 wpscbe2 = 5.899567621e-15 ppscbe2 = -1.756743748e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.467571504e-08 lalpha0 = 3.548251731e-14 walpha0 = 3.197479574e-13 palpha0 = -1.751499374e-19   alpha1 = 5.130872968e-10 lalpha1 = -2.262788940e-16 walpha1 = -2.039094733e-15 palpha1 = 1.116965117e-21   beta0 = -2.341150040e+01 lbeta0 = 1.768417239e-05 wbeta0 = 1.626828886e-04 pbeta0 = -8.836203145e-11   agidl = 1.0e-10   bgidl = 9.772225167e+08 lbgidl = 1.112143628e+02 wbgidl = 7.263893590e+02 pbgidl = -4.402227599e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.202537151e-01 lkt1 = -3.713388333e-08 wkt1 = -4.326050283e-07 pkt1 = 2.281071748e-13   kt2 = -2.273752259e-02 lkt2 = -3.324924039e-09 wkt2 = -2.171375431e-08 pkt2 = -2.762991932e-15   at = -4.732749015e+04 lat = 3.343866352e-02 wat = 5.620443105e-01 pat = -2.080118330e-7   ute = -1.138512217e-01 lute = 2.109602991e-09 wute = -4.689917886e-07 pute = 2.569019770e-13   ua1 = 4.576679483e-09 lua1 = -1.024469240e-15 wua1 = -2.678541710e-15 pua1 = 9.355286546e-22   ub1 = -4.973910940e-18 lub1 = 1.367407035e-24 wub1 = 8.962320017e-24 pub1 = -3.414546503e-30   uc1 = -3.484286942e-10 luc1 = 6.577897655e-17 wuc1 = 6.070022280e-17 puc1 = 9.219306096e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.213288245e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.578202867e-08 wvth0 = 6.658240729e-07 pvth0 = -1.633462660e-13   k1 = -8.807755003e-01 lk1 = 4.750807296e-07 wk1 = 5.944787091e-06 pk1 = -1.703022895e-12   k2 = 5.187223371e-01 lk2 = -1.754422763e-07 wk2 = -2.052780889e-06 pk2 = 5.873278470e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 4.160470621e+00 ldsub = -1.063508820e-06 wdsub = -2.144186162e-05 pdsub = 6.580170386e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.139655356e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.545204206e-08 wvoff = -2.630893559e-07 pvoff = 4.565341897e-14   nfactor = {6.693685792e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.189892084e-06 wnfactor = -2.996178054e-05 pnfactor = 7.270479275e-12   eta0 = 0.49   etab = -6.249996614e-04 letab = -1.008117418e-16 wetab = -1.671161598e-15 petab = 4.976301454e-22   u0 = 1.859294642e-02 lu0 = -4.267118927e-09 wu0 = -7.821666609e-08 pu0 = 2.415334169e-14   ua = 2.715906428e-09 lua = -1.417615811e-15 wua = -2.281960518e-14 pua = 7.224357254e-21   ub = -1.915118612e-18 lub = 1.108324938e-24 wub = 1.641115777e-23 pub = -5.144790732e-30   uc = 7.381768986e-11 luc = -1.200098990e-17 wuc = -2.645049267e-16 puc = 9.580975727e-24   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.482549449e+05 lvsat = -4.679870429e-02 wvsat = -1.381694679e+00 pvsat = 3.847576762e-7   a0 = 4.113985297e+00 la0 = -9.644600525e-07 wa0 = -1.911687923e-05 pa0 = 5.500140126e-12   ags = 9.346321080e+00 lags = -1.844139534e-06 wags = -2.499347544e-05 pags = 5.692888869e-12   a1 = 0.0   a2 = -1.981574403e-01 la2 = 2.972263318e-07 wa2 = 8.625496167e-06 pa2 = -2.568457121e-12   b0 = 0.0   b1 = 0.0   keta = 4.322488014e-01 lketa = -1.453010977e-07 wketa = -3.588908640e-06 pketa = 1.003023322e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.265258665e+00 lpclm = -9.967429308e-08 wpclm = -3.338944022e-06 ppclm = 5.639033676e-13   pdiblc1 = 9.701137241e-01 lpdiblc1 = -1.379196406e-07 wpdiblc1 = -4.868723499e-06 ppdiblc1 = 1.176870579e-12   pdiblc2 = 4.693323123e-03 lpdiblc2 = 1.080812381e-09 wpdiblc2 = 1.117126675e-08 ppdiblc2 = -3.021378018e-15   pdiblcb = 1.032062508e+00 lpdiblcb = -3.147667882e-07 wpdiblcb = -3.937721873e-06 ppdiblcb = 1.172555131e-12   drout = 4.006117051e-01 ldrout = 1.347744730e-07 wdrout = 6.028678342e-07 pdrout = -7.806959406e-13   pscbe1 = 7.983276287e+08 lpscbe1 = 4.979903646e-01 wpscbe1 = 1.390796390e+01 ppscbe1 = -4.141443951e-6   pscbe2 = -7.313237347e-08 lpscbe2 = 2.207476751e-14 wpscbe2 = 3.272700605e-13 ppscbe2 = -9.745284227e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 6.880390652e-08 lalpha0 = -4.264377003e-15 walpha0 = -3.391384219e-13 palpha0 = 2.104995422e-20   alpha1 = -2.468116000e-10 walpha1 = 1.711942518e-15   beta0 = 4.367681487e+01 lbeta0 = -2.293050692e-06 wbeta0 = -1.769947542e-04 pbeta0 = 1.278547864e-11   agidl = 1.0e-10   bgidl = -1.549775331e+09 lbgidl = 8.636911469e+02 wbgidl = 1.586889863e+04 pbgidl = -4.949283459e-3   cgidl = 3.132084150e+03 lcgidl = -8.433238577e-04 wcgidl = -1.397982441e-02 pcgidl = 4.162842213e-9   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.927548560e-01 lkt1 = -4.532235607e-08 wkt1 = -2.527585662e-07 pkt1 = 1.745533945e-13   kt2 = 2.851534031e-02 lkt2 = -1.858674529e-08 wkt2 = -1.318400732e-07 pkt2 = 3.002987267e-14   at = 1.287413118e+05 lat = -1.899022398e-02 wat = -3.021743296e-01 pat = 4.933087257e-8   ute = -1.812805381e+00 lute = 5.080156778e-07 wute = 1.486656330e-05 pute = -4.309642940e-12   ua1 = 3.604876788e-09 lua1 = -7.350906927e-16 wua1 = 1.970369958e-15 pua1 = -4.488010172e-22   ub1 = -1.853443330e-18 lub1 = 4.382097923e-25 wub1 = -1.065416657e-23 pub1 = 2.426752790e-30   uc1 = -5.120450788e-10 luc1 = 1.144998455e-16 wuc1 = 1.575258140e-15 puc1 = -3.588044229e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-6.999859201e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.719095410e-08 wvth0 = -1.948243555e-06 pvth0 = 4.643207798e-13   k1 = 2.343450373e+00 lk1 = -2.786714814e-07 wk1 = -1.430313362e-05 pk1 = 3.126056686e-12   k2 = -1.964660237e-01 lk2 = -1.347618948e-08 wk2 = 3.102615286e-06 pk2 = -6.307490048e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -6.579123681e+00 ldsub = 1.485900335e-06 wdsub = 6.225311860e-05 pdsub = -1.341515701e-11   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.334478079e-03+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.467614876e-08 wvoff = -9.880686573e-07 pvoff = 2.265175730e-13   nfactor = {-1.460956394e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.935803206e-06 wnfactor = 8.501118568e-05 pnfactor = -2.032939590e-11   eta0 = 2.421684939e+00 leta0 = -4.728281808e-07 weta0 = 8.948165329e-09 peta0 = -2.190287168e-15   etab = 4.175968295e-01 letab = -1.023702483e-07 wetab = -1.151488051e-06 petab = 2.818554879e-13   u0 = -6.098314964e-02 lu0 = 1.489264333e-08 wu0 = 3.805855884e-07 pu0 = -8.634729414e-14   ua = -2.074955754e-08 lua = 4.220339295e-15 wua = 1.086414980e-13 pua = -2.441484397e-20   ub = 1.442276598e-17 lub = -2.808060869e-24 wub = -7.074753852e-23 pub = 1.580549740e-29   uc = 3.635087585e-10 luc = -8.380581579e-17 wuc = -2.395195977e-15 puc = 5.318359543e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.944962250e+04 lvsat = 1.523585726e-02 wvsat = 2.356894427e+00 pvsat = -5.016390612e-7   a0 = -9.151029076e-01 la0 = 1.945524821e-07 wa0 = 1.113635185e-05 pa0 = -1.494591244e-12   ags = 1.25   a1 = 0.0   a2 = 3.536357312e+00 la2 = -5.947060126e-07 wa2 = -2.244524300e-05 pa2 = 4.845186115e-12   b0 = -5.232177336e-23 lb0 = 1.280706207e-29 wb0 = 2.582724120e-28 pb0 = -6.321862964e-35   b1 = 0.0   keta = -1.283430862e+00 lketa = 2.638098363e-07 wketa = 4.987061297e-06 pketa = -1.021299017e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.237646620e+00 lpclm = -3.451297511e-07 wpclm = -6.901772797e-06 ppclm = 1.478081741e-12   pdiblc1 = 1.214372709e+00 lpdiblc1 = -2.080017739e-07 wpdiblc1 = 5.774804345e-06 ppdiblc1 = -1.340563146e-12   pdiblc2 = 4.091813931e-02 lpdiblc2 = -7.705450507e-09 wpdiblc2 = 4.175716148e-08 ppdiblc2 = -1.073354112e-14   pdiblcb = -3.137311828e+00 lpdiblcb = 6.822991779e-07 wpdiblcb = 2.021483495e-05 ppdiblcb = -4.651873247e-12   drout = 9.372701190e-01 ldrout = 1.347281020e-08 wdrout = -2.304654174e-05 pdrout = 4.949821002e-12   pscbe1 = 8.041934406e+08 lpscbe1 = -9.006462053e-01 wpscbe1 = -3.487396634e+01 ppscbe1 = 7.490056120e-6   pscbe2 = 1.238015403e-07 lpscbe2 = -2.448217971e-14 wpscbe2 = -8.058865170e-13 ppscbe2 = 1.726421606e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.705078021e-07 lalpha0 = -5.395472006e-14 walpha0 = -1.334795646e-12 palpha0 = 2.663330157e-19   alpha1 = -2.468116000e-10 walpha1 = 1.711942518e-15   beta0 = 7.352237738e+01 lbeta0 = -9.769640224e-06 wbeta0 = -2.816402119e-04 pbeta0 = 3.935431545e-11   agidl = 1.0e-10   bgidl = 5.442474586e+09 lbgidl = -7.833751889e+02 wbgidl = -2.244482102e+04 pbgidl = 4.059567217e-3   cgidl = -6.801399458e+03 lcgidl = 1.525203069e-03 wcgidl = 3.505415525e-02 pcgidl = -7.528756193e-9   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -9.003151537e-01 lkt1 = 7.553307917e-08 wkt1 = 3.192762239e-06 pkt1 = -6.557961581e-13   kt2 = -1.012651270e+00 lkt2 = 2.348775890e-07 wkt2 = 6.034649561e-06 pkt2 = -1.477131346e-12   at = 5.409557811e+05 lat = -1.213073572e-01 wat = -3.114074941e+00 pat = 7.412956572e-7   ute = 6.616547734e+00 lute = -1.517363452e-06 wute = -4.143755181e-05 pute = 9.150546392e-12   ua1 = -3.847987056e-09 lua1 = 1.034320519e-15 wua1 = 2.755779995e-14 pua1 = -6.745460482e-21   ub1 = 6.307372079e-18 lub1 = -1.526647987e-24 wub1 = -3.769590826e-23 pub1 = 9.227015944e-30   uc1 = 6.553525337e-10 luc1 = -1.627042027e-16 wuc1 = -3.257789106e-15 puc1 = 7.974253284e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.094192049e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.303952113e-08 wvth0 = -6.807168019e-09 pvth0 = 6.810420144e-13   k1 = 4.561927827e-01 lk1 = -1.963033664e-06 wk1 = -9.389344432e-08 pk1 = 9.393830191e-12   k2 = 3.041826054e-02 lk2 = 8.411822293e-07 wk2 = 4.193453405e-08 pk2 = -4.195456827e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.635402555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.786910346e-07 wvoff = -1.175911352e-08 pvoff = 1.176473144e-12   nfactor = {2.045336893e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.467126075e-05 wnfactor = -1.944390916e-06 pnfactor = 1.945319848e-10   eta0 = 0.08   etab = -0.07   u0 = 9.167404527e-03 lu0 = 1.802795603e-08 wu0 = 1.154371695e-09 pu0 = -1.154923196e-13   ua = -1.037912001e-10 lua = 5.123869774e-15 wua = 3.175539068e-16 pua = -3.177056182e-20   ub = 1.250771594e-19 lub = -4.838853595e-24 wub = -2.851716694e-25 pub = 2.853079102e-29   uc = -8.810478989e-11 luc = 1.043907878e-15 wuc = 5.383830284e-17 puc = -5.386402409e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.099455759e+05 lvsat = -9.950327378e-1   a0 = 1.534471683e+00 la0 = 6.354466119e-06 wa0 = 1.501920999e-07 pa0 = -1.502638542e-11   ags = 2.317150564e-01 lags = 3.393494831e-06 wags = -2.312110743e-08 pags = 2.313215354e-12   a1 = 0.0   a2 = 1.050106932e+00 la2 = -5.014087489e-6   b0 = 0.0   b1 = 0.0   keta = 3.020738088e-03 lketa = -1.619755477e-06 wketa = -3.424324052e-08 pketa = 3.425960023e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 8.012853566e-03 lpclm = 6.750904548e-06 wpclm = 2.094174854e-07 ppclm = -2.095175346e-11   pdiblc1 = 0.39   pdiblc2 = 4.539339641e-03 lpdiblc2 = -9.121758245e-08 wpdiblc2 = -2.190217888e-10 ppdiblc2 = 2.191264264e-14   pdiblcb = 1.213132527e-03 lpdiblcb = -1.309501882e-07 wpdiblcb = -2.787585881e-09 ppdiblcb = 2.788917651e-13   drout = 0.56   pscbe1 = 7.797360482e+08 lpscbe1 = -3.327680857e+03 wpscbe1 = -1.298788880e+02 ppscbe1 = 1.299409376e-2   pscbe2 = 9.390041541e-09 lpscbe2 = 1.150058773e-14 wpscbe2 = 4.438158047e-16 ppscbe2 = -4.440278377e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.316586945e-10 lalpha0 = 2.317693695e-14 walpha0 = 6.802036719e-16 palpha0 = -6.805286392e-20   alpha1 = 1.616800379e-10 lalpha1 = -6.170950555e-15 walpha1 = -1.811069011e-16 palpha1 = 1.811934249e-20   beta0 = 5.108713286e+00 lbeta0 = -3.164753098e-05 wbeta0 = 3.900592812e-07 pbeta0 = -3.902456320e-11   agidl = 1.168985839e-10 lagidl = -1.690665723e-15 wagidl = -8.341533075e-17 pagidl = 8.345518242e-21   bgidl = 9.145685115e+08 lbgidl = 2.399906893e+04 wbgidl = 8.179739569e+02 pbgidl = -8.183647439e-2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.529705238e-01 lkt1 = 1.128591306e-06 wkt1 = 4.331322393e-08 pkt1 = -4.333391682e-12   kt2 = -0.037961   at = 0.0   ute = -2.803718620e-01 lute = -2.029783062e-06 wute = -3.821007260e-08 pute = 3.822832746e-12   ua1 = 2.317372900e-09 lua1 = -1.058234334e-14 wua1 = -5.221195757e-16 pua1 = 5.223690183e-20   ub1 = -1.041468335e-18 lub1 = 2.479967592e-23 wub1 = 1.380647604e-24 pub1 = -1.381307209e-28   uc1 = 2.324401938e-10 luc1 = -1.126439837e-14 wuc1 = -5.557713174e-16 puc1 = 5.560368371e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.098832939e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.716378459e-8   k1 = 3.582750006e-01 wk1 = 3.746787634e-7   k2 = 7.237714272e-02 wk2 = -1.673384066e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.874177698e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = 4.692436351e-8   nfactor = {-1.829034361e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 7.759029282e-6   eta0 = 0.08   etab = -0.07   u0 = 1.006665425e-02 wu0 = -4.606483043e-9   ua = 1.517917648e-10 wua = -1.267188631e-15   ub = -1.162889571e-19 wub = 1.137968356e-24   uc = -3.603378061e-11 wuc = -2.148400123e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160312.5   a0 = 1.851437836e+00 wa0 = -5.993367340e-7   ags = 4.009854533e-01 wags = 9.226403402e-8   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -7.777403727e-02 wketa = 1.366465476e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 3.447536913e-01 wpclm = -8.356737261e-7   pdiblc1 = 0.39   pdiblc2 = -1.067064477e-05 wpdiblc2 = 8.739993890e-10   pdiblcb = -5.318773791e-03 wpdiblcb = 1.112377162e-8   drout = 0.56   pscbe1 = 6.137485080e+08 wpscbe1 = 5.182775166e+2   pscbe2 = 9.963700599e-09 wpscbe2 = -1.771032664e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.024426554e-09 walpha0 = -2.714330830e-15   alpha1 = -1.461322034e-10 walpha1 = 7.227012517e-16   beta0 = 3.530107631e+00 wbeta0 = -1.556518990e-6   agidl = 3.256674547e-11 wagidl = 3.328661889e-16   bgidl = 2.111662400e+09 wbgidl = -3.264098712e+3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.966754334e-01 wkt1 = -1.728400241e-7   kt2 = -0.037961   at = 0.0   ute = -3.816191606e-01 wute = 1.524760632e-7   ua1 = 1.789516650e-09 wua1 = 2.083501339e-15   ub1 = 1.955605078e-19 wub1 = -5.509429767e-24   uc1 = -3.294375395e-10 wuc1 = 2.217787530e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.094554632e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.443085161e-08 wvth0 = -2.848367630e-08 pvth0 = 4.478382446e-13   k1 = 2.609826751e-01 lk1 = 7.829867448e-07 wk1 = 5.602878804e-07 pk1 = -1.493740412e-12   k2 = 1.176093365e-01 lk2 = -3.640185185e-07 wk2 = -2.767513015e-07 pk2 = 8.805303602e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.689287847e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.487951921e-07 wvoff = -2.642261417e-08 pvoff = 5.902799733e-13   nfactor = {2.007924158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.087897885e-06 wnfactor = 7.378823089e-06 pnfactor = 3.059813891e-12   eta0 = 0.08   etab = -0.07   u0 = 8.367301161e-03 lu0 = 1.367601127e-08 wu0 = 7.379060116e-09 pu0 = -9.645695460e-14   ua = -3.363994309e-10 lua = 3.928852899e-15 wua = 2.118336272e-15 pua = -2.724594268e-20   ub = 2.118396561e-19 lub = -2.640705250e-24 wub = -1.025812917e-24 pub = 1.741362483e-29   uc = 4.368331852e-11 luc = -6.415452775e-16 wuc = -5.476169325e-16 puc = 2.678113779e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.315729531e+05 lvsat = -5.734880933e-01 wvsat = -2.764463862e-02 pvsat = 2.224778316e-7   a0 = 1.501998120e+00 la0 = 2.812212211e-06 wa0 = 5.361564486e-07 pa0 = -9.138193648e-12   ags = 4.016274341e-02 lags = 2.903819984e-06 wags = 1.153323118e-06 pags = -8.539164773e-12   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -6.479969098e-02 lketa = -1.044146196e-07 wketa = 8.007834902e-08 pketa = 4.552481347e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.325438018e-02 lpclm = 2.345920868e-06 wpclm = -1.681328530e-06 ppclm = 6.805639592e-12   pdiblc1 = 0.39   pdiblc2 = -2.390366433e-04 lpdiblc2 = 1.837838174e-09 wpdiblc2 = 1.758437608e-09 ppdiblc2 = -7.117759790e-15   pdiblcb = -6.970151752e-03 lpdiblcb = 1.328991828e-08 wpdiblcb = 1.920361045e-08 ppdiblcb = -6.502472500e-14   drout = 0.56   pscbe1 = 6.150978036e+08 lpscbe1 = -1.085882691e+01 wpscbe1 = 4.853740055e+02 ppscbe1 = 2.648000536e-4   pscbe2 = 1.165112574e-08 lpscbe2 = -1.358001785e-14 wpscbe2 = -7.344052427e-15 ppscbe2 = 4.485040912e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.959894228e-09 lalpha0 = -7.528433358e-15 walpha0 = -5.461080948e-15 palpha0 = 2.210522694e-20   alpha1 = -3.952041482e-10 lalpha1 = 2.004474971e-15 walpha1 = 1.454034267e-15 palpha1 = -5.885603553e-21   beta0 = 2.137801120e+00 lbeta0 = 1.120496953e-05 wbeta0 = -8.439114231e-06 pbeta0 = 5.538957791e-11   agidl = -9.387504891e-09 lagidl = 7.581061702e-14 wagidl = 2.812885929e-14 pagidl = -2.236958984e-19   bgidl = 9.661008581e+08 lbgidl = 9.219221537e+03 wbgidl = -4.896561326e+02 pbgidl = -2.232808963e-2   cgidl = 300.0   egidl = -4.239518307e-01 legidl = 4.216646444e-06 wegidl = 1.538444132e-06 pegidl = -1.238105222e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.054705530e-01 lkt1 = -7.339963563e-07 wkt1 = -6.033174762e-07 pkt1 = 3.464385677e-12   kt2 = -3.129229069e-02 lkt2 = -5.366827209e-8   at = -1.906940243e+05 lat = 1.534662601e+00 wat = 2.684067248e-02 pat = -2.160076930e-7   ute = 9.874183524e-01 lute = -1.101770587e-05 wute = -2.403107966e-06 pute = 2.056676526e-11   ua1 = 3.942231319e-09 lua1 = -1.732456329e-14 wua1 = 4.191887497e-15 pua1 = -1.696781741e-20   ub1 = -1.712235121e-19 lub1 = 2.951795266e-24 wub1 = -1.201169268e-23 pub1 = 5.232874890e-29   uc1 = -7.241740676e-10 luc1 = 3.176750762e-15 wuc1 = 4.462063759e-15 puc1 = -1.806143013e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.139254685e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.465049024e-07 wvth0 = 2.822775286e-07 pvth0 = -8.100531916e-13   k1 = 2.344075660e-01 lk1 = 8.905568071e-07 wk1 = 1.073675313e-06 pk1 = -3.571817226e-12   k2 = 9.987499185e-02 lk2 = -2.922338815e-07 wk2 = -3.220218715e-07 pk2 = 1.063775442e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.469062737e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.668401385e-07 wvoff = 3.402677505e-07 pvoff = -8.940001176e-13   nfactor = {-2.252234145e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.841401703e-06 wnfactor = 1.573190247e-05 pnfactor = -3.075157201e-11   eta0 = 0.08   etab = -0.07   u0 = 1.987441571e-02 lu0 = -3.290219933e-08 wu0 = -5.013330575e-08 pu0 = 1.363401621e-13   ua = 2.637764325e-09 lua = -8.109892798e-15 wua = -1.191941118e-14 pua = 2.957570054e-20   ub = -1.515607075e-18 lub = 4.351610440e-24 wub = 6.347240066e-24 pub = -1.243083471e-29   uc = -2.087178439e-10 luc = 3.801178379e-16 wuc = 4.170496918e-16 puc = -1.226639666e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.722338118e+05 lvsat = -3.332966006e-01 wvsat = -7.688448246e-02 pvsat = 4.217896405e-7   a0 = 1.817651064e+00 la0 = 1.534520113e-06 wa0 = 7.353136981e-07 pa0 = -9.944337384e-12   ags = 6.057523495e-02 lags = 2.821194811e-06 wags = 1.360152078e-06 pags = -9.376361863e-12   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -3.550009684e-02 lketa = -2.230127843e-07 wketa = -1.809152813e-08 pketa = 8.526177091e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.236974266e-01 lpclm = 3.689576620e-08 wpclm = 9.361693845e-07 ppclm = -3.789403030e-12   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = -4.114443565e-02 lpdiblcb = 1.516197303e-07 wpdiblcb = 1.804127695e-07 ppdiblcb = -7.175631289e-13   drout = 0.56   pscbe1 = 4.216893736e+08 lpscbe1 = 7.720149809e+02 wpscbe1 = 1.110807767e+03 ppscbe1 = -2.266815092e-3   pscbe2 = -2.538213451e-09 lpscbe2 = 4.385523459e-14 wpscbe2 = 5.716527788e-14 ppscbe2 = -2.162688454e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -2.801102260e-03 lalpha0 = 1.133823210e-08 walpha0 = 8.224686384e-09 palpha0 = -3.329167993e-14   alpha1 = 3.527073121e-10 lalpha1 = -1.022902340e-15 walpha1 = -7.420072964e-16 palpha1 = 3.003478584e-21   beta0 = -6.492801546e+01 lbeta0 = 2.826723052e-04 wbeta0 = 2.068886844e-04 pbeta0 = -8.162089020e-10   agidl = 1.880366595e-08 lagidl = -3.830089955e-14 wagidl = -5.491830249e-14 pagidl = 1.124603269e-19   bgidl = 5.078131610e+09 lbgidl = -7.425353738e+03 wbgidl = -1.155922633e+04 pbgidl = 2.247903989e-2   cgidl = 300.0   egidl = 1.147903661e+00 legidl = -2.145870920e-06 wegidl = -3.076888263e-06 pegidl = 6.300774864e-12   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.562846892e-01 lkt1 = 2.812428338e-07 wkt1 = 6.298158862e-07 pkt1 = -1.527060719e-12   kt2 = -3.965545262e-02 lkt2 = -1.981607430e-08 wkt2 = -1.140732337e-09 pkt2 = 4.617427836e-15   at = 3.731235917e+05 lat = -7.475442492e-01 wat = -2.810179931e-01 pat = 1.030134917e-6   ute = -3.339788572e+00 lute = 6.497854135e-06 wute = 4.918721762e-06 pute = -9.070354069e-12   ua1 = -2.403186070e-09 lua1 = 8.360258579e-15 wua1 = -2.813890526e-15 pua1 = 1.138999572e-20   ub1 = 2.142939302e-18 lub1 = -6.415415119e-24 wub1 = 3.216163322e-24 pub1 = -9.310185919e-30   uc1 = 2.818507105e-11 luc1 = 1.313702500e-16 wuc1 = 1.905998149e-16 puc1 = -7.715051658e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.026734937e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.391022379e-08 wvth0 = -2.711551928e-07 pvth0 = 3.232524996e-13   k1 = 9.210155439e-01 lk1 = -5.154618448e-07 wk1 = -1.436500138e-06 pk1 = 1.568457308e-12   k2 = -1.208872985e-01 lk2 = 1.598376177e-07 wk2 = 4.375638703e-07 pk2 = -4.916852505e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 6.320709603e-02 ldsub = 1.017320089e-06 wdsub = 9.349886265e-07 pdsub = -1.914646335e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.375584702e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.707955982e-08 wvoff = -2.149040900e-07 pvoff = 2.428668981e-13   nfactor = {6.373941377e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.240931460e-07 wnfactor = 9.102540706e-07 pnfactor = -4.001709551e-13   eta0 = -6.823364663e-02 leta0 = 3.035491557e-07 weta0 = 7.627202217e-09 peta0 = -1.561879402e-14   etab = -6.390916566e-01 letab = 1.165371667e-06 wetab = 4.017691184e-06 petab = -8.227327564e-12   u0 = -3.867842821e-03 lu0 = 1.571660414e-08 wu0 = 4.210603178e-08 pu0 = -5.254524727e-14   ua = -2.373576705e-09 lua = 2.152206080e-15 wua = 6.575842275e-15 pua = -8.298417116e-21   ub = 4.896207774e-19 lub = 2.453549758e-25 wub = -1.052766518e-25 pub = 7.824677144e-31   uc = 2.506646473e-11 luc = -9.861982480e-17 wuc = -4.365510550e-16 puc = 5.213426034e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.611989787e+04 lvsat = 1.547981673e-01 wvsat = 3.104305577e-01 pvsat = -3.713444158e-7   a0 = 4.048682252e+00 la0 = -3.034129777e-06 wa0 = -8.604021444e-06 pa0 = 9.180519637e-12   ags = 2.382963083e+00 lags = -1.934532965e-06 wags = -6.714899265e-06 pags = 7.159526401e-12   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -2.835599545e-01 lketa = 2.849579907e-07 wketa = 8.259502137e-07 pketa = -8.757898687e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 7.098524234e-01 lpclm = -1.395302824e-07 wpclm = -2.014252658e-06 ppclm = 2.252397469e-12   pdiblc1 = 3.769517587e-01 lpdiblc1 = 2.671986239e-08 wpdiblc1 = 9.681629469e-08 ppdiblc1 = -1.982579879e-13   pdiblc2 = -1.027162500e-05 lpdiblc2 = 4.613056019e-10   pdiblcb = 9.355955857e-02 lpdiblcb = -1.242237415e-07 wpdiblcb = -3.481183698e-07 ppdiblcb = 3.647497249e-13   drout = 8.532238145e-01 ldrout = -6.004563968e-07 wdrout = -2.185051974e-06 pdrout = 4.474494806e-12   pscbe1 = 7.973199379e+08 lpscbe1 = 2.808102096e+00 wpscbe1 = 7.869284181e+00 ppscbe1 = -8.245239233e-6   pscbe2 = 2.912798146e-08 lpscbe2 = -2.099000769e-14 wpscbe2 = -9.979997434e-14 ppscbe2 = 1.051606740e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 5.565623084e-03 lalpha0 = -5.794938887e-09 walpha0 = -1.634196031e-08 palpha0 = 1.701528500e-14   alpha1 = -1.468116000e-10 walpha1 = 7.246961179e-16   beta0 = 9.073361548e+01 lbeta0 = -3.608769106e-05 wbeta0 = -2.466453731e-04 pbeta0 = 1.125268025e-10   agidl = 1.0e-10   bgidl = 1.259250660e+09 lbgidl = 3.948551992e+02 wbgidl = 3.154574436e+01 pbgidl = -1.256253401e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.430147935e-01 lkt1 = -1.554859268e-07 wkt1 = -2.954273560e-07 pkt1 = 3.676292612e-13   kt2 = -3.807881310e-02 lkt2 = -2.304467730e-08 wkt2 = -6.756064865e-08 pkt2 = 1.406304720e-13   at = -1.074828201e+05 lat = 2.366295457e-01 wat = 5.029659512e-01 pat = -5.752878045e-7   ute = 3.367085960e+00 lute = -7.236315859e-06 wute = -9.886545542e-06 pute = 2.124750219e-11   ua1 = 8.143133554e-09 lua1 = -1.323623109e-14 wua1 = -1.558066734e-14 pua1 = 3.753348211e-20   ub1 = -4.948473762e-18 lub1 = 8.106203269e-24 wub1 = 1.003135619e-23 pub1 = -2.326616750e-29   uc1 = -4.599627213e-11 luc1 = 2.832769501e-16 wuc1 = 6.055271352e-16 puc1 = -1.621182959e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.114060851e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.587686380e-09 wvth0 = -3.650223072e-08 pvth0 = 7.738899217e-14   k1 = 5.074294416e-01 lk1 = -8.211666645e-08 wk1 = -5.539138552e-07 pk1 = 6.437054653e-13   k2 = 1.409351624e-03 lk2 = 3.169824511e-08 wk2 = 1.878694552e-07 pk2 = -2.300616848e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.071543808e+00 ldsub = -3.918990939e-08 wdsub = -1.869977253e-06 pdsub = 1.024326790e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.457663567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.847954163e-08 wvoff = -1.235021507e-07 pvoff = 1.470982312e-13   nfactor = {3.158649853e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.717615561e-06 wnfactor = -4.032047525e-06 pnfactor = 4.778249099e-12   eta0 = 4.389143691e-01 leta0 = -2.278278565e-07 weta0 = -1.875722198e-07 peta0 = 1.889062803e-13   etab = 9.910289442e-01 letab = -5.426279454e-07 wetab = -8.032406751e-06 petab = 4.398463800e-12   u0 = 1.252891616e-02 lu0 = -1.463510008e-09 wu0 = -5.136950539e-09 pu0 = -3.045231470e-15   ua = 1.001931184e-09 lua = -1.384566698e-15 wua = -3.828071184e-15 pua = 2.602543309e-21   ub = -1.003909170e-18 lub = 1.810238316e-24 wub = 5.130972133e-24 pub = -4.703942856e-30   uc = -1.670752004e-10 luc = 1.027014084e-16 wuc = 2.963572338e-16 puc = -2.465803789e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -5.735474518e+03 lvsat = 9.152887813e-02 wvsat = 1.903021927e-01 pvsat = -2.454769182e-7   a0 = 8.836310719e-01 la0 = 2.821317233e-07 wa0 = 1.032725833e-06 pa0 = -9.166232407e-13   ags = 1.629373259e-01 lags = 3.915545230e-07 wags = -9.591444185e-07 pags = 1.128790366e-12   a1 = 0.0   a2 = 1.037062068e+00 la2 = -2.483877085e-07 wa2 = -1.339394856e-06 pa2 = 1.403384446e-12   b0 = 0.0   b1 = 0.0   keta = -1.264281314e-02 lketa = 1.097782900e-09 wketa = 9.608450513e-08 pketa = -1.110548259e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.439106514e-01 lpclm = -7.043814219e-08 wpclm = -3.413691863e-07 ppclm = 4.995919886e-13   pdiblc1 = 1.380229911e+00 lpdiblc1 = -1.024489904e-06 wpdiblc1 = -4.986793284e-06 ppdiblc1 = 5.128221039e-12   pdiblc2 = -1.804765749e-03 lpdiblc2 = 2.341531682e-09 wpdiblc2 = 4.671741577e-09 ppdiblc2 = -4.894934031e-15   pdiblcb = 1.467303428e-02 lpdiblcb = -4.156841350e-08 wpdiblcb = -1.958353014e-07 ppdiblcb = 2.051913329e-13   drout = 2.392875695e-01 ldrout = 4.281065233e-08 wdrout = 2.267018200e-06 pdrout = -1.902730200e-13   pscbe1 = 7.859334965e+08 lpscbe1 = 1.473853067e+01 wpscbe1 = 6.943552455e+01 ppscbe1 = -7.275280674e-5   pscbe2 = 8.789795948e-09 lpscbe2 = 3.198346298e-16 wpscbe2 = 1.623428112e-15 ppscbe2 = -1.108231497e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 7.316357109e-05 lalpha0 = -4.007712037e-11 walpha0 = -2.148249250e-10 palpha0 = 1.176757233e-16   alpha1 = -4.172060484e-10 lalpha1 = 2.833125432e-16 walpha1 = 1.518636950e-15 palpha1 = -8.318713552e-22   beta0 = 1.081489569e+02 lbeta0 = -5.433505045e-05 wbeta0 = -2.928501212e-04 pbeta0 = 1.609389825e-10   agidl = 1.0e-10   bgidl = 2.202600608e+09 lbgidl = -5.935632925e+02 wbgidl = -2.692934830e+03 pbgidl = 1.598389233e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.916664990e-01 lkt1 = 2.676139275e-10 wkt1 = 1.169543444e-07 pkt1 = -6.445397491e-14   kt2 = -1.098957583e-01 lkt2 = 5.220332244e-08 wkt2 = 2.458572672e-07 pkt2 = -1.877609848e-13   at = 1.673651904e+05 lat = -5.134932859e-02 wat = 2.765849078e-02 pat = -7.727253018e-8   ute = -7.151468730e+00 lute = 3.784762782e-06 wute = 2.106270711e-05 pute = -1.118035101e-11   ua1 = -1.273433947e-08 lua1 = 8.638663212e-15 wua1 = 4.526317467e-14 pua1 = -2.621717444e-20   ub1 = 8.355375679e-18 lub1 = -5.833237580e-24 wub1 = -2.750550590e-23 pub1 = 1.606401818e-29   uc1 = 8.491940819e-10 luc1 = -6.546811231e-16 wuc1 = -2.860445180e-15 puc1 = 2.010376184e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.144424027e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.421987472e-08 wvth0 = 2.664943768e-07 pvth0 = -8.858497449e-14   k1 = -2.709561557e-01 lk1 = 3.442635041e-07 wk1 = 2.094881038e-06 pk1 = -8.072381572e-13   k2 = 2.914440633e-01 lk2 = -1.271755191e-07 wk2 = -7.961194516e-07 pk2 = 3.089428386e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.093869945e+00 ldsub = -5.141960901e-08 wdsub = 1.172128889e-06 pdsub = -6.420629022e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.308904488e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.850692056e-09 wvoff = 2.270809766e-07 pvoff = -4.494244138e-14   nfactor = {-9.805786494e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.497503319e-07 wnfactor = 6.111860711e-06 pnfactor = -7.783302345e-13   eta0 = -5.332451517e-01 leta0 = 3.046968251e-07 weta0 = 3.446356306e-07 peta0 = -1.026238749e-13   etab = 1.676175446e-03 letab = -6.852325185e-10 wetab = -5.951233280e-09 petab = 1.772128490e-15   u0 = 1.806193379e-02 lu0 = -4.494358740e-09 wu0 = -3.449494087e-08 pu0 = 1.303634169e-14   ua = -6.544456103e-10 lua = -4.772448996e-16 wua = -9.430945152e-16 pua = 1.022225214e-21   ub = 2.907361447e-18 lub = -3.322579456e-25 wub = -6.631677757e-24 pub = 1.739342687e-30   uc = 5.041576887e-11 luc = -1.643470732e-17 wuc = -2.853813661e-16 puc = 7.208148263e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.795343076e+05 lvsat = -6.473477675e-02 wvsat = -6.284687209e-01 pvsat = 2.030253190e-7   a0 = 2.233637850e+00 la0 = -4.573682396e-07 wa0 = -1.677230890e-06 pa0 = 5.678233033e-13   ags = 1.084785861e-01 lags = 4.213856592e-07 wags = -1.699342101e-07 pags = 6.964807442e-13   a1 = 0.0   a2 = 3.258758636e-01 la2 = 1.411823147e-07 wa2 = 2.678789713e-06 pa2 = -7.976766066e-13   b0 = 0.0   b1 = 0.0   keta = 1.541384030e-01 lketa = -9.026079776e-08 wketa = -5.194288558e-07 pketa = 2.261080054e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 3.709568459e-01 lpclm = 7.907912857e-08 wpclm = 1.243181497e-06 ppclm = -3.683852620e-13   pdiblc1 = -1.358450379e+00 lpdiblc1 = 4.756906923e-07 wpdiblc1 = 9.102767868e-06 ppdiblc1 = -2.589688321e-12   pdiblc2 = -5.648106796e-03 lpdiblc2 = 4.446817825e-09 wpdiblc2 = -4.905444017e-09 ppdiblc2 = 3.512088080e-16   pdiblcb = -1.043460686e-01 lpdiblcb = 2.362727557e-08 wpdiblcb = 3.916706027e-07 ppdiblcb = -1.166297137e-13   drout = 1.562591464e-01 ldrout = 8.829154683e-08 wdrout = 4.256395258e-06 pdrout = -1.280004038e-12   pscbe1 = 8.278753575e+08 lpscbe1 = -8.236172200e+00 wpscbe1 = -1.375992315e+02 ppscbe1 = 4.065565677e-5   pscbe2 = 3.358318669e-08 lpscbe2 = -1.326136499e-14 wpscbe2 = -7.114618660e-14 ppscbe2 = 3.875314420e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.944357401e+00 lbeta0 = 6.749057178e-09 wbeta0 = 2.966867879e-06 pbeta0 = -1.102168721e-12   agidl = 1.0e-10   bgidl = 7.472986600e+08 lbgidl = 2.036147319e+02 wbgidl = 1.861346858e+03 pbgidl = -8.963324185e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.277408549e-01 lkt1 = 2.002824419e-08 wkt1 = 9.797643081e-08 pkt1 = -5.405834827e-14   kt2 = -1.119881765e-03 lkt2 = -7.381383316e-09 wkt2 = -1.284234447e-07 pkt2 = 1.726063216e-14   at = 1.283442596e+05 lat = -2.997463820e-02 wat = -3.051122022e-01 pat = 1.050109362e-7   ute = -4.511581370e-01 lute = 1.145001467e-07 wute = 1.196033400e-06 pute = -2.978838214e-13   ua1 = 6.149374868e-09 lua1 = -1.705363412e-15 wua1 = -1.044173099e-14 pua1 = 4.296580254e-21   ub1 = -4.936420944e-18 lub1 = 1.447676316e-24 wub1 = 8.777260703e-24 pub1 = -3.810774297e-30   uc1 = -8.089355198e-10 luc1 = 2.536008195e-16 wuc1 = 2.333868752e-15 puc1 = -8.349391303e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.018143727e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.338324164e-08 wvth0 = -2.974545412e-07 pvth0 = 7.934491457e-14   k1 = 1.173592627e+00 lk1 = -8.588700973e-08 wk1 = -4.196050599e-06 pk1 = 1.066044011e-12   k2 = -2.150098627e-01 lk2 = 2.363379872e-08 wk2 = 1.569091475e-06 pk2 = -3.953578450e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -1.426189704e+00 ldsub = 6.989911528e-07 wdsub = 6.135189844e-06 pdsub = -2.119938378e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.799454999e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.702082420e-08 wvoff = 6.260305550e-08 pvoff = 4.034971571e-15   nfactor = {-7.134223254e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.701978575e-07 wnfactor = 6.601423571e-06 pnfactor = -9.241098151e-13   eta0 = 0.49   etab = -0.000625   u0 = -1.016836641e-02 lu0 = 3.911918904e-09 wu0 = 6.375584670e-08 pu0 = -1.622028658e-14   ua = -5.008657242e-09 lua = 8.193304691e-16 wua = 1.531063320e-14 pua = -3.817728555e-21   ub = 2.582808942e-18 lub = -2.356143236e-25 wub = -5.791656159e-24 pub = 1.489205256e-30   uc = 1.321257106e-10 luc = -4.076588522e-17 wuc = -5.523268446e-16 puc = 1.515711725e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.206259691e+05 lvsat = 5.442294963e-02 wvsat = 4.391870929e-01 pvsat = -1.148958910e-7   a0 = -6.287910605e-01 la0 = 3.949915292e-07 wa0 = 4.294565190e-06 pa0 = -1.210428274e-12   ags = 2.413844574e+00 lags = -2.650946979e-07 wags = 9.226836926e-06 pags = -2.101642781e-12   a1 = 0.0   a2 = 1.994111536e+00 la2 = -3.555765627e-07 wa2 = -2.196052108e-06 pa2 = 6.539294164e-13   b0 = 0.0   b1 = 0.0   keta = -6.564317070e-01 lketa = 1.511067167e-07 wketa = 1.785070924e-06 pketa = -4.601144165e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.749206564e-01 lpclm = -1.007661951e-07 wpclm = -1.905768251e-06 ppclm = 5.692932492e-13   pdiblc1 = -1.914955573e-01 lpdiblc1 = 1.282007202e-07 wpdiblc1 = 8.652494068e-07 ppdiblc1 = -1.367612617e-13   pdiblc2 = 1.430017107e-02 lpdiblc2 = -1.493280618e-09 wpdiblc2 = -3.625036353e-08 ppdiblc2 = 9.684942215e-15   pdiblcb = -3.385040258e-01 lpdiblcb = 9.335366128e-08 wpdiblcb = 2.827712507e-06 ppdiblcb = -8.420220917e-13   drout = 1.821792396e+00 ldrout = -4.076626165e-07 wdrout = -6.412409769e-06 pdrout = 1.896899379e-12   pscbe1 = 8.037465523e+08 lpscbe1 = -1.051217236e+00 wpscbe1 = -1.284110008e+01 ppscbe1 = 3.505804180e-6   pscbe2 = -2.942803358e-08 lpscbe2 = 5.501801133e-15 wpscbe2 = 1.115352994e-13 ppscbe2 = -1.564483530e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.601109903e+00 lbeta0 = 4.067345810e-07 wbeta0 = 1.083295057e-06 pbeta0 = -5.412878235e-13   agidl = 1.153599337e-09 lagidl = -3.137355425e-16 wagidl = -5.200810761e-15 pagidl = 1.548671424e-21   bgidl = 2.392420652e+09 lbgidl = -2.862614693e+02 wbgidl = -3.590695327e+03 pbgidl = 7.271494431e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.066134079e-01 lkt1 = 1.373701867e-08 wkt1 = 3.092736610e-07 pkt1 = -1.169773810e-13   kt2 = 8.303888093e-02 lkt2 = -3.244175888e-08 wkt2 = -4.009809191e-07 pkt2 = 9.842143410e-14   at = -6.018439496e+04 lat = 2.616448191e-02 wat = 6.304067897e-01 pat = -1.735632316e-7   ute = 2.863524793e+00 lute = -8.725295627e-07 wute = -8.216887346e-06 pute = 2.505048654e-12   ua1 = 2.840773108e-09 lua1 = -7.201445229e-16 wua1 = 5.742162997e-15 pua1 = -5.225787789e-22   ub1 = -3.124901682e-18 lub1 = 9.082511672e-25 wub1 = -4.377953168e-24 pub1 = 1.065195138e-31   uc1 = 1.314066773e-10 luc1 = -2.640957828e-17 wuc1 = -1.600969009e-15 puc1 = 3.367571839e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.146680850e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.708057365e-08 wvth0 = 2.567462507e-07 pvth0 = -5.038767211e-14   k1 = -1.474257289e+00 lk1 = 5.558302716e-07 wk1 = 4.541957111e-06 pk1 = -9.932375713e-13   k2 = 8.052505124e-01 lk2 = -2.243365247e-07 wk2 = -1.842089935e-06 pk2 = 4.101065294e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.121999155e+01 ldsub = -2.344308620e-06 wdsub = -2.560744360e-05 pdsub = 5.491643002e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.504344090e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.551475166e-08 wvoff = -2.570130389e-07 pvoff = 8.257015141e-14   nfactor = {-6.180847628e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.819548493e-07 wnfactor = 1.594599845e-05 pnfactor = -3.280399118e-12   eta0 = 2.424068936e+00 leta0 = -4.734117237e-07 weta0 = -2.819797728e-09 peta0 = 6.902159889e-16   etab = 4.577587234e-01 letab = -1.122008759e-07 wetab = -1.349736477e-06 petab = 3.303817462e-13   u0 = 2.598873459e-02 lu0 = -4.646469205e-09 wu0 = -4.872780960e-08 pu0 = 1.010229838e-14   ua = 3.502563119e-09 lua = -1.202852719e-15 wua = -1.107259603e-14 pua = 2.355289993e-21   ub = -8.850892852e-19 lub = 5.956553767e-25 wub = 4.815586489e-24 pub = -9.960356447e-31   uc = -3.037713355e-10 luc = 6.288825009e-17 wuc = 8.986533758e-16 puc = -1.922799879e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.461056743e+05 lvsat = -1.047144285e-01 wvsat = -4.348177275e-01 pvsat = 9.046337765e-8   a0 = 3.691838958e+00 la0 = -6.331104684e-07 wa0 = -1.160458201e-05 pa0 = 2.590945097e-12   ags = 1.25   a1 = 0.0   a2 = -2.435744082e+00 la2 = 7.022028694e-07 wa2 = 7.034435013e-06 pa2 = -1.556657010e-12   b0 = 0.0   b1 = 0.0   keta = 8.913526776e-02 lketa = -2.011158116e-08 wketa = -1.788243554e-06 pketa = 3.802029693e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.213802367e-01 lpclm = 1.600601654e-07 wpclm = 4.742931061e-06 ppclm = -1.015652891e-12   pdiblc1 = 2.040456517e+00 lpdiblc1 = -4.085570808e-07 wpdiblc1 = 1.697063017e-06 ppdiblc1 = -3.505756226e-13   pdiblc2 = 4.034316826e-02 lpdiblc2 = -7.979406338e-09 wpdiblc2 = 4.459535194e-08 ppdiblc2 = -9.381231578e-15   pdiblcb = -6.917344157e+00 lpdiblcb = 1.710656710e-06 wpdiblcb = 3.887395150e-05 ppdiblcb = -9.728084606e-12   drout = -6.897810176e+00 ldrout = 1.696252180e-06 wdrout = 1.562923233e-05 pdrout = -3.356768374e-12   pscbe1 = 7.929129147e+08 lpscbe1 = 1.522128751e+00 wpscbe1 = 2.080932672e+01 ppscbe1 = -4.469323146e-6   pscbe2 = -1.112784588e-07 lpscbe2 = 2.594736621e-14 wpscbe2 = 3.545228972e-13 ppscbe2 = -7.628977771e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.797500458e+01 lbeta0 = -2.102178829e-06 wbeta0 = -7.445492698e-06 pbeta0 = 1.505947152e-12   agidl = -2.215923311e-09 lagidl = 4.876236938e-16 wagidl = 1.143193476e-14 pagidl = -2.407023681e-21   bgidl = 7.421320966e+08 lbgidl = 9.632277091e+01 wbgidl = 7.571599899e+02 pbgidl = -2.828260023e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.048153947e-01 lkt1 = -8.358782685e-08 wkt1 = -7.340091273e-07 pkt1 = 1.296615501e-13   kt2 = 5.439061853e-01 lkt2 = -1.476718458e-07 wkt2 = -1.648879161e-06 pkt2 = 4.112214156e-13   at = -1.186104293e+05 lat = 4.241850206e-02 wat = 1.416968933e-01 pat = -6.689316835e-8   ute = -7.081222424e+00 lute = 1.496574644e-06 wute = 2.617781958e-05 pute = -5.726951285e-12   ua1 = -1.547610480e-09 lua1 = 3.002740427e-16 wua1 = 1.620260748e-14 pua1 = -3.122036775e-21   ub1 = 8.492719249e-19 lub1 = 3.260199884e-27 wub1 = -1.075345962e-23 pub1 = 1.675034195e-30   uc1 = 2.788144945e-11 luc1 = -3.040271006e-18 wuc1 = -1.604462608e-16 puc1 = 9.287119644e-24   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.100849615e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.258966318e-07 wvth0 = 1.274099114e-08 pvth0 = -2.554285237e-13   k1 = 4.300098230e-01 lk1 = 1.120078752e-06 wk1 = -1.701420013e-08 pk1 = 3.410968559e-13   k2 = 4.554497998e-02 lk2 = -6.046149116e-07 wk2 = -2.481023628e-09 pk2 = 4.973900346e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.443312138e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.434030846e-07 wvoff = -6.816131645e-08 pvoff = 1.366482736e-12   nfactor = {1.891364221e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.139204146e-05 wnfactor = -1.492291432e-06 pnfactor = 2.991712286e-11   eta0 = 0.08   etab = -0.07   u0 = 1.007908518e-02 lu0 = -3.170099697e-08 wu0 = -1.522534222e-09 pu0 = 3.052342351e-14   ua = 1.311046807e-10 lua = -8.237281328e-15 wua = -3.721548951e-16 pua = 7.460877602e-21   ub = -6.292891566e-20 lub = 6.699981153e-24 wub = 2.668577843e-25 pub = -5.349904817e-30   uc = -6.520169976e-11 luc = -8.821159378e-16 wuc = -1.341048330e-17 puc = 2.688503519e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.060467257e+05 lvsat = -2.921646966e+00 wvsat = -2.821752712e-01 pvsat = 5.656986348e-6   a0 = 1.265904905e+00 la0 = 7.646528007e-06 wa0 = 9.387664657e-07 pa0 = -1.882017888e-11   ags = -1.491658220e-01 lags = 1.165926213e-05 wags = 1.095233516e-06 pags = -2.195699510e-11   a1 = 0.0   a2 = 1.534371976e+00 la2 = -1.472252414e-05 wa2 = -1.421914519e-06 pa2 = 2.850622235e-11   b0 = 0.0   b1 = 0.0   keta = 8.076451381e-02 lketa = -2.245360599e-06 wketa = -2.625170026e-07 pketa = 5.262881801e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.627377178e-01 lpclm = 4.468325933e-06 wpclm = 7.107807771e-07 ppclm = -1.424957309e-11   pdiblc1 = 0.39   pdiblc2 = 1.284588590e-02 lpdiblc2 = -2.517779282e-07 wpdiblc2 = -2.460896872e-08 ppdiblc2 = 4.933550679e-13   pdiblcb = 7.454327465e-03 lpdiblcb = -1.801222430e-07 wpdiblcb = -2.111318218e-08 ppdiblcb = 4.232723258e-13   drout = 0.56   pscbe1 = 8.026545589e+08 lpscbe1 = -2.484913464e+02 wpscbe1 = -1.971729525e+02 ppscbe1 = 3.952878987e-3   pscbe2 = 9.299228060e-09 lpscbe2 = 1.229077765e-15 wpscbe2 = 7.104652527e-16 ppscbe2 = -1.424324753e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -8.069465346e-10 lalpha0 = 1.818226006e-14 walpha0 = 2.663005437e-15 palpha0 = -5.338733383e-20   alpha1 = 3.414780795e-10 lalpha1 = -4.841098204e-15 walpha1 = -7.090356642e-16 palpha1 = 1.421458746e-20   beta0 = 9.061646906e+00 lbeta0 = -1.215225333e-04 wbeta0 = -1.121667091e-05 pbeta0 = 2.248692946e-10   agidl = 8.848961259e-11 lagidl = 1.151588650e-15   bgidl = 4.764853565e+08 lbgidl = 1.049530378e+04 wbgidl = 2.104287735e+03 pbgidl = -4.218628705e-2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.624336919e-01 lkt1 = 1.382031839e-07 wkt1 = 7.109928093e-08 pkt1 = -1.425382387e-12   kt2 = -0.037961   at = 0.0   ute = -1.721433477e-01 lute = -3.158459837e-06 wute = -3.559940996e-07 pute = 7.136889611e-12   ua1 = 2.139553309e-09 lua1 = 7.208111171e-15   ub1 = -2.638066334e-19 lub1 = -2.840756419e-23 wub1 = -9.027475700e-25 pub1 = 1.809808017e-29   uc1 = 4.315974271e-11 luc1 = 7.672689606e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.0895817+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.4858803   k2 = 0.015386276   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.17143662+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.4596089+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.0084978126   ua = -2.7977789e-10   ub = 2.7127182e-19   uc = -1.0920239e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160312.5   a0 = 1.6473202   ags = 0.43240805   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -0.031235975   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.060146165   pdiblc1 = 0.39   pdiblc2 = 0.00028698955   pdiblcb = -0.0015303226   drout = 0.56   pscbe1 = 790259600.0   pscbe2 = 9.3605355e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   agidl = 1.4593183e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.45554   kt2 = -0.037961   at = 0.0   ute = -0.32969   ua1 = 2.4991e-9   ub1 = -1.6808e-18   uc1 = 4.2588e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.104255390e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.180905583e-7   k1 = 4.518013436e-01 lk1 = 2.742597737e-7   k2 = 2.335544192e-02 lk2 = -6.413405423e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.779276016e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.223795970e-8   nfactor = {2.713816962e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.045809286e-6   eta0 = 0.08   etab = -0.07   u0 = 1.088040643e-02 lu0 = -1.917457908e-8   ua = 3.850477410e-10 lua = -5.350367093e-15   ub = -1.375240580e-19 lub = 3.289897247e-24   uc = -1.428199730e-10 luc = 2.705467437e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.221579483e+05 lvsat = -4.977182523e-1   a0 = 1.684598285e+00 la0 = -3.000056410e-7   ags = 4.329529311e-01 lags = -4.385080593e-9   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -3.752720400e-02 lketa = 5.063039543e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.193599535e-01 lpclm = 4.663734853e-06 ppclm = 8.881784197e-28   pdiblc1 = 0.39   pdiblc2 = 3.598389252e-04 lpdiblc2 = -5.862753804e-10   pdiblcb = -4.299292994e-04 lpdiblcb = -8.855717695e-9   drout = 0.56   pscbe1 = 7.804028631e+08 lpscbe1 = 7.932480083e+1   pscbe2 = 9.149943124e-09 lpscbe2 = 1.694800055e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -7.363294768e-01 lbeta0 = 3.006913896e-5   agidl = 1.924122583e-10 lagidl = -3.740640288e-16   bgidl = 7.993374236e+08 lbgidl = 1.614887265e+3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.109439203e-01 lkt1 = 4.458782848e-7   kt2 = -3.129229069e-02 lkt2 = -5.366827209e-8   at = -1.815528282e+05 lat = 1.461096312e+0   ute = 1.689857606e-01 lute = -4.013230319e-6   ua1 = 5.369873105e-09 lua1 = -2.310333602e-14   ub1 = -4.262076237e-18 lub1 = 2.077353037e-23 pub1 = -1.232595164e-44   uc1 = 7.954823353e-10 luc1 = -2.974476434e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.043118709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.293769733e-7   k1 = 6.000718980e-01 lk1 = -3.259060697e-7   k2 = -9.796815934e-03 lk2 = 7.005882629e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.310204205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.376317553e-7   nfactor = {3.105619891e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.631739389e-6   eta0 = 0.08   etab = -0.07   u0 = 2.800388268e-03 lu0 = 1.353151645e-8   ua = -1.421659857e-09 lua = 1.962778754e-15 wua = 1.654361225e-30   ub = 6.460886178e-19 lub = 1.180094484e-25   uc = -6.668216971e-11 luc = -3.764195286e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.460490681e+05 lvsat = -1.896466300e-1   a0 = 2.068078721e+00 la0 = -1.852248161e-6   ags = 5.238056873e-01 lags = -3.721365957e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -4.166157459e-02 lketa = 6.736539737e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.425310148e-01 lpclm = -1.253670861e-6   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = 2.029920012e-02 lpdiblcb = -9.276256952e-08 wpdiblcb = 3.469446952e-24 ppdiblcb = -4.163336342e-29   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.693071063e-08 lpscbe2 = -2.979999612e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.532589957e+00 lbeta0 = 4.693963595e-6   agidl = 1.0e-10   bgidl = 1.141376499e+09 lbgidl = 2.303900486e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.417866910e-01 lkt1 = -2.388321190e-7   kt2 = -4.004395473e-02 lkt2 = -1.824350515e-8   at = 2.774165791e+05 lat = -3.967085806e-1   ute = -1.664606991e+00 lute = 3.408740581e-6   ua1 = -3.361519923e-09 lua1 = 1.223937839e-14 wua1 = 8.271806126e-31 pua1 = 4.963083675e-36   ub1 = 3.238276224e-18 lub1 = -9.586208816e-24 pub1 = -3.081487911e-45   uc1 = 9.309813477e-11 luc1 = -1.313832265e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.119082951e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.618070211e-8   k1 = 4.317830385e-01 lk1 = 1.871164947e-8   k2 = 2.813494163e-02 lk2 = -7.616878557e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 3.816385505e-01 ldsub = 3.652441172e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.107489027e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.563423735e-8   nfactor = {9.474016816e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.878059061e-7   eta0 = -6.563603097e-02 leta0 = 2.982298233e-07 peta0 = -1.110223025e-28   etab = 7.292236481e-01 letab = -1.636630206e-06 wetab = -2.220446049e-22   u0 = 1.047231551e-02 lu0 = -2.178864366e-9   ua = -1.340253773e-10 lua = -6.740069421e-16   ub = 4.537664404e-19 lub = 5.118419953e-25   uc = -1.236108384e-10 luc = 7.893515158e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.960422667e+04 lvsat = 2.832845517e-2   a0 = 1.118388786e+00 la0 = 9.250314490e-8   ags = 9.605276213e-02 lags = 5.038051506e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -2.263989568e-03 lketa = -1.331199231e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.385327269e-02 lpclm = 6.275744520e-7   pdiblc1 = 4.099247304e-01 lpdiblc1 = -4.080136477e-8   pdiblc2 = -1.027162500e-05 lpdiblc2 = 4.613056019e-10   pdiblcb = -0.025   drout = 1.090551064e-01 ldrout = 9.234336795e-7   pscbe1 = 800000000.0   pscbe2 = -4.861149626e-09 lpscbe2 = 1.482483051e-14 ppscbe2 = -3.308722450e-36   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.732973460e+00 lbeta0 = 2.235848267e-6   agidl = 1.0e-10   bgidl = 1.269994274e+09 lbgidl = -3.299021648e+1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.436292395e-01 lkt1 = -3.028149435e-8   kt2 = -6.108811503e-02 lkt2 = 2.485020020e-8   at = 6.381357310e+04 lat = 4.070231495e-2   ute = 0.0   ua1 = 2.836786052e-09 lua1 = -4.533576282e-16   ub1 = -1.532069271e-18 lub1 = 1.823854303e-25   uc1 = 1.602296443e-10 luc1 = -2.688534535e-16 wuc1 = 5.169878828e-32 puc1 = 5.169878828e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.126492509e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.394425227e-8   k1 = 3.187815911e-01 lk1 = 1.371117410e-7   k2 = 6.539252981e-02 lk2 = -4.665444801e-08 pk2 = 2.775557562e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 4.346808990e-01 ldsub = 3.096676706e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.878277982e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.618077084e-9   nfactor = {1.785445172e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.027511255e-8   eta0 = 3.750324212e-01 leta0 = -1.634915641e-7   etab = -1.744588252e+00 letab = 9.553680575e-7   u0 = 1.077941185e-02 lu0 = -2.500632234e-9   ua = -3.018047553e-10 lua = -4.982119042e-16   ub = 7.435590590e-19 lub = 2.082045343e-25   uc = -6.614406353e-11 luc = 1.872290159e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.907622725e+04 lvsat = 7.926179768e-3   a0 = 1.235349135e+00 la0 = -3.004498506e-8   ags = -1.637209281e-01 lags = 7.759895289e-07 pags = -4.440892099e-28   a1 = 0.0   a2 = 5.809009555e-01 la2 = 2.295665014e-7   b0 = 0.0   b1 = 0.0   keta = 2.008093115e-02 lketa = -3.672444161e-08 pketa = -1.387778781e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.276496794e-01 lpclm = 9.970917197e-8   pdiblc1 = -3.181349608e-01 lpdiblc1 = 7.220413781e-7   pdiblc2 = -2.136988382e-04 lpdiblc2 = 6.744515502e-10   pdiblcb = -5.202309237e-02 lpdiblcb = 2.831412061e-8   drout = 1.011371724e+00 ldrout = -2.199111402e-8   pscbe1 = 8.095813297e+08 lpscbe1 = -1.003907775e+1   pscbe2 = 9.342690989e-09 lpscbe2 = -5.759858989e-17   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.412246329e+00 lbeta0 = 4.763481371e-7   agidl = 1.0e-10   bgidl = 1.285460944e+09 lbgidl = -4.919580623e+1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.518350605e-01 lkt1 = -2.168364023e-8   kt2 = -2.616352350e-02 lkt2 = -1.174291369e-8   at = 1.767849130e+05 lat = -7.766623072e-2   ute = 2.191100000e-02 lute = -2.295779803e-8   ua1 = 2.681055040e-09 lua1 = -2.901865670e-16   ub1 = -1.012244420e-18 lub1 = -3.622740528e-25   uc1 = -1.249950081e-10 luc1 = 2.999780679e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.053663359e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.949735344e-9   k1 = 4.425028073e-01 lk1 = 6.934035184e-8   k2 = 2.030763693e-02 lk2 = -2.195807082e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.493064862e+00 ldsub = -2.700886046e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.535529031e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.715685362e-8   nfactor = {1.100953297e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.846724244e-7   eta0 = -4.158717185e-01 leta0 = 2.697459510e-07 weta0 = -1.110223025e-22 peta0 = -1.110223025e-28   etab = -3.506512077e-04 letab = -8.169421162e-11   u0 = 6.313904049e-03 lu0 = -5.453869694e-11   ua = -9.756377079e-10 lua = -1.291030586e-16   ub = 6.487940866e-19 lub = 2.601144171e-25   uc = -4.677728878e-11 luc = 8.114266548e-18 wuc = -5.169878828e-32   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.549511688e+04 lvsat = 4.410072501e-3   a0 = 1.662419060e+00 la0 = -2.639832131e-7   ags = 5.060366000e-02 lags = 6.585878776e-7   a1 = 0.0   a2 = 1.238198089e+00 la2 = -1.304844360e-7   b0 = 0.0   b1 = 0.0   keta = -2.276480350e-02 lketa = -1.325461931e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 7.943503302e-01 lpclm = -4.638277703e-8   pdiblc1 = 1.741702425e+00 lpdiblc1 = -4.062860457e-07 ppdiblc1 = 4.440892099e-28   pdiblc2 = -7.318766341e-03 lpdiblc2 = 4.566429902e-09 wpdiblc2 = -3.469446952e-24 ppdiblc2 = -4.336808690e-31   pdiblcb = 2.904618475e-02 lpdiblcb = -1.609360266e-08 wpdiblcb = 6.938893904e-24 ppdiblcb = -6.505213035e-31   drout = 1.605870505e+00 ldrout = -3.476426838e-07 wdrout = -1.776356839e-21   pscbe1 = 7.810128372e+08 lpscbe1 = 5.610028227e+0   pscbe2 = 9.352748976e-09 lpscbe2 = -6.310810356e-17   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.954791140e+00 lbeta0 = -3.686193471e-7   agidl = 1.0e-10   bgidl = 1.381222293e+09 lbgidl = -1.016514795e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.943727726e-01 lkt1 = 1.617455029e-9   kt2 = -4.485738095e-02 lkt2 = -1.502885923e-9   at = 2.443142092e+04 lat = 5.789203407e-3   ute = -4.382200000e-02 lute = 1.304909605e-8   ua1 = 2.593207986e-09 lua1 = -2.420661471e-16   ub1 = -1.947126944e-18 lub1 = 1.498312215e-25   uc1 = -1.408390333e-11 luc1 = -3.075652365e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.119448738e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.363950580e-08 wvth0 = 4.741177868e-13 pvth0 = -1.411804238e-19   k1 = -2.554668373e-01 lk1 = 2.771782628e-07 wk1 = -4.697547631e-13 pk1 = 1.398812239e-19   k2 = 3.193795685e-01 lk2 = -1.110142152e-07 wk2 = 1.263829361e-13 pk2 = -3.763367873e-20   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 6.632874742e-01 ldsub = -2.300164303e-08 wdsub = 9.176943117e-14 pdsub = -2.732664228e-20   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.586246647e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.564660981e-08 wvoff = 1.367088132e-13 pvoff = -4.070846660e-20   nfactor = {1.534841430e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.554713858e-07 wnfactor = -4.112898466e-13 pnfactor = 1.224718336e-19   eta0 = 0.49   etab = -0.000625   u0 = 1.154512665e-02 lu0 = -1.612266006e-09 wu0 = -6.457309909e-15 pu0 = 1.922825461e-21   ua = 2.057241424e-10 lua = -4.808830836e-16 wua = -2.850525139e-22 pua = 8.488151079e-29   ub = 6.103299983e-19 lub = 2.715680610e-25 wub = -3.638200364e-31 pub = 1.083365114e-37   uc = -5.598164756e-11 luc = 1.085509448e-17 wuc = -8.726124737e-26 puc = 2.598425043e-32   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.894910005e+04 lvsat = 1.529256266e-02 wvsat = -1.148423017e-08 pvsat = 3.419716610e-15   a0 = 8.338199239e-01 la0 = -1.724710534e-08 wa0 = 1.367088487e-14 pa0 = -4.070847659e-21   ags = 5.556251721e+00 lags = -9.808564737e-07 wags = 5.046590559e-13 pags = -1.502748503e-19   a1 = 0.0   a2 = 1.246196109e+00 la2 = -1.328660465e-07 wa2 = 1.101814867e-12 pa2 = -3.280929208e-19   b0 = 0.0   b1 = 0.0   keta = -4.848556225e-02 lketa = -5.595620375e-09 wketa = -7.271752089e-16 pketa = 2.165346236e-22   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 3.258683178e-01 lpclm = 9.311945420e-08 wpclm = -4.799353803e-15 ppclm = 1.429127039e-21   pdiblc1 = 1.031846539e-01 lpdiblc1 = 8.162358351e-08 wpdiblc1 = -5.890113464e-14 ppdiblc1 = 1.753928514e-20   pdiblc2 = 1.954292813e-03 lpdiblc2 = 1.805144712e-09 wpdiblc2 = -7.068137187e-16 ppdiblc2 = 2.104714528e-22   pdiblcb = 6.245371022e-01 lpdiblcb = -1.934159106e-07 wpdiblcb = 3.295554976e-13 ppdiblcb = -9.813338800e-20   drout = -3.620983483e-01 ldrout = 2.383692413e-07 wdrout = 1.183840119e-13 pdrout = -3.525179970e-20   pscbe1 = 7.993732294e+08 lpscbe1 = 1.427624370e-01 wpscbe1 = -9.598705292e-06 ppscbe1 = 2.858254433e-12   pscbe2 = 8.557826678e-09 lpscbe2 = 1.735998837e-16 wpscbe2 = 9.845943007e-22 ppscbe2 = -2.931875705e-28   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.970050275e+00 lbeta0 = 2.223868641e-07 wbeta0 = 5.308374398e-13 pbeta0 = -1.580701223e-19   agidl = -6.176539417e-10 lagidl = 2.136994025e-16 wagidl = -2.050632297e-22 pagidl = 6.106270309e-29   bgidl = 1.169528257e+09 lbgidl = -3.861428793e+01 wbgidl = 4.552112617e-04 pbgidl = -1.355505333e-10   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.012832461e-01 lkt1 = -2.610227873e-08 wkt1 = -1.306005419e-13 pkt1 = 3.888957645e-20   kt2 = -5.352420734e-02 lkt2 = 1.077878303e-09 wkt2 = -9.358735786e-15 pkt2 = 2.786797570e-21   at = 1.545148243e+05 lat = -3.294638204e-02 wat = 7.169941068e-08 pat = -2.135029199e-14   ute = 6.507857669e-02 lute = -1.937877317e-08 wute = -1.544518813e-14 pute = 4.599190903e-21   ua1 = 4.796396516e-09 lua1 = -8.981206116e-16 wua1 = -1.034042205e-21 pua1 = 3.079119148e-28   ub1 = -4.615912639e-18 lub1 = 9.445288819e-25 wub1 = 9.162399519e-31 pub1 = -2.728333511e-37   uc1 = -4.138393819e-10 luc1 = 8.828066398e-17 wuc1 = -8.217072412e-23 puc1 = 2.446838726e-29   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.059240368e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.001267327e-11 wvth0 = 7.098486776e-13 pvth0 = -2.094184630e-19   k1 = 7.260845696e-02 lk1 = 2.175608479e-07 wk1 = 4.088205330e-13 pk1 = -6.473200109e-20   k2 = 1.778849916e-01 lk2 = -8.466543241e-08 wk2 = 7.833103952e-13 pk2 = -2.012418894e-19   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.498799548e+00 ldsub = -4.740058399e-07 wdsub = -5.531242273e-13 pdsub = 1.284876774e-19   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.379658463e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.606342309e-09 wvoff = -4.319228033e-13 pvoff = 9.544005852e-20   nfactor = {4.812683932e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.352588972e-07 wnfactor = 1.617939617e-12 pnfactor = -3.650921165e-19   eta0 = 2.423108485e+00 leta0 = -4.731766295e-07 weta0 = 3.078033757e-13 peta0 = -7.534257218e-20   etab = -1.924461846e-03 letab = 3.180757735e-10 wetab = 1.055179354e-15 petab = -2.582815264e-22   u0 = 9.393374142e-03 lu0 = -1.205902351e-09 wu0 = 1.879193604e-14 pu0 = -4.114048539e-21   ua = -2.684595089e-10 lua = -4.007055165e-16 wua = 1.281320490e-21 pua = -2.921923035e-28   ub = 7.549669653e-19 lub = 2.564330450e-25 wub = 8.439094927e-31 pub = -1.791997849e-37   uc = 2.285327712e-12 luc = -2.597033798e-18 wuc = 7.553276462e-24 puc = -1.842289073e-30   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.980184987e+05 lvsat = -7.390503813e-02 wvsat = 5.762362313e-07 pvsat = -1.401843285e-13   a0 = -2.603633681e-01 la0 = 2.492943713e-07 wa0 = 9.339082112e-13 pa0 = -2.296257664e-19   ags = 1.250000431e+00 lags = -9.256125200e-14 wags = -1.265423400e-12 pags = 2.717813086e-19   a1 = 0.0   a2 = -4.000781802e-02 la2 = 1.720480550e-07 wa2 = -2.469248098e-12 pa2 = 5.215267800e-19   b0 = 0.0   b1 = 0.0   keta = -5.198915673e-01 lketa = 1.093751551e-07 wketa = 5.279603341e-13 pketa = -1.291767894e-19   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.493931515e+00 lpclm = -1.858432392e-07 wpclm = 1.005943460e-12 ppclm = -2.458687822e-19   pdiblc1 = 2.618430104e+00 lpdiblc1 = -5.279536407e-07 wpdiblc1 = -1.523348889e-12 ppdiblc1 = 3.773085293e-19   pdiblc2 = 5.553109607e-02 lpdiblc2 = -1.117439023e-08 wpdiblc2 = 7.230731697e-14 ppdiblc2 = -1.764585383e-20   pdiblcb = 6.322061588e+00 lpdiblcb = -1.602463074e-06 wpdiblcb = -1.531498873e-11 ppdiblcb = 3.723935734e-18   drout = -1.574923469e+00 ldrout = 5.530292122e-07 wdrout = 2.054833470e-12 pdrout = -5.118772357e-19   pscbe1 = 7.999999918e+08 lpscbe1 = 1.760531425e-06 wpscbe1 = 2.406857300e-05 ppscbe1 = -5.169328690e-12   pscbe2 = 9.462306747e-09 lpscbe2 = -3.483758818e-17 wpscbe2 = -2.389380683e-21 ppscbe2 = 5.107950661e-28   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.543927404e+01 lbeta0 = -1.589294526e-06 wbeta0 = 4.489302796e-13 pbeta0 = -1.498188595e-19   agidl = 1.677480134e-09 lagidl = -3.321425738e-16 wagidl = -1.024909967e-21 pagidl = 2.662981068e-28   bgidl = 1.000000389e+09 lbgidl = -8.349186230e-05 wbgidl = -1.141433960e-03 pbgidl = 2.451514778e-10   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.547988797e-01 lkt1 = -3.942863456e-08 wkt1 = 3.808868847e-13 pkt1 = -8.340723401e-20   kt2 = -1.765682813e-02 lkt2 = -7.621111934e-09 wkt2 = 1.290873346e-13 pkt2 = -3.089334666e-20   at = -7.035235195e+04 lat = 1.963652595e-02 wat = -1.776520442e-08 pat = -1.045071098e-15   ute = 1.834224364e+00 lute = -4.538677692e-07 wute = -5.808090946e-13 pute = 1.433294021e-19   ua1 = 3.970551439e-09 lua1 = -7.630056656e-16 wua1 = 3.872934809e-21 pua1 = -8.702123579e-28   ub1 = -2.813060016e-18 lub1 = 5.737305977e-25 wub1 = -3.378441247e-30 pub1 = 7.580343072e-37   uc1 = -2.676221162e-11 luc1 = 1.226819692e-19 wuc1 = 2.054006927e-22 puc1 = -4.409570666e-29   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.094269313e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.397621949e-8   k1 = 4.212225495e-01 lk1 = 1.296244034e-6   k2 = 4.426361306e-02 lk2 = -5.789263560e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.795342868e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.623402023e-7   nfactor = {1.120644890e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.684324920e-5   eta0 = 0.08   etab = -0.07   u0 = 9.292746448e-03 lu0 = -1.593665493e-08 wu0 = 1.387778781e-23   ua = -6.110105453e-11 lua = -4.383983995e-15 pua = -3.308722450e-36   ub = 7.489433296e-20 lub = 3.936931675e-24   uc = -7.212777231e-11 luc = -7.432635937e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160312.5   a0 = 1.750746838e+00 la0 = -2.073473977e-6   ags = 4.164861845e-01 lags = 3.191979779e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -5.481686414e-02 lketa = 4.727443598e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.043571226e-01 lpclm = -2.891108831e-6   pdiblc1 = 0.39   pdiblc2 = 1.361647904e-04 lpdiblc2 = 3.023700845e-9   pdiblcb = -3.449935132e-03 lpdiblcb = 3.848396013e-8   drout = 0.56   pscbe1 = 7.008212287e+08 lpscbe1 = 1.793040344e+3   pscbe2 = 9.666159942e-09 lpscbe2 = -6.127090055e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 5.684079876e-10 lalpha0 = -9.390537943e-15   alpha1 = -2.471546770e-11 lalpha1 = 2.500267635e-15 walpha1 = -2.019483917e-33 palpha1 = 3.231174268e-37   beta0 = 3.268606140e+00 lbeta0 = -5.384955464e-6   agidl = 8.848961259e-11 lagidl = 1.151588650e-15   bgidl = 1.563280604e+09 lbgidl = -1.129252281e+4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.257132571e-01 lkt1 = -5.979598311e-7   kt2 = -0.037961   at = 0.0   ute = -3.560025648e-01 lute = 5.275083793e-7   ua1 = 2.139553309e-09 lua1 = 7.208111171e-15   ub1 = -7.300459942e-19 lub1 = -1.906050239e-23 wub1 = 1.540743956e-39   uc1 = 4.315974271e-11 luc1 = 7.672689606e-15 puc1 = -6.617444900e-36   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.0895817+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.4858803   k2 = 0.015386276   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.17143662+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.4596089+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.0084978126   ua = -2.7977789e-10   ub = 2.7127182e-19   uc = -1.0920239e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160312.5   a0 = 1.6473202   ags = 0.43240805   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -0.031235975   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.060146165   pdiblc1 = 0.39   pdiblc2 = 0.00028698955   pdiblcb = -0.0015303226   drout = 0.56   pscbe1 = 790259600.0   pscbe2 = 9.3605355e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   agidl = 1.4593183e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.45554   kt2 = -0.037961   at = 0.0   ute = -0.32969   ua1 = 2.4991e-9   ub1 = -1.6808e-18   uc1 = 4.2588e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.104255390e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.180905583e-7   k1 = 4.518013436e-01 lk1 = 2.742597737e-7   k2 = 2.335544192e-02 lk2 = -6.413405423e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.779276016e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.223795970e-8   nfactor = {2.713816962e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.045809286e-6   eta0 = 0.08   etab = -0.07   u0 = 1.088040643e-02 lu0 = -1.917457908e-8   ua = 3.850477410e-10 lua = -5.350367093e-15   ub = -1.375240580e-19 lub = 3.289897247e-24 pub = 3.081487911e-45   uc = -1.428199730e-10 luc = 2.705467437e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.221579483e+05 lvsat = -4.977182523e-01 wvsat = 4.656612873e-16   a0 = 1.684598285e+00 la0 = -3.000056410e-7   ags = 4.329529311e-01 lags = -4.385080593e-9   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -3.752720400e-02 lketa = 5.063039543e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.193599535e-01 lpclm = 4.663734853e-06 wpclm = 2.220446049e-22 ppclm = -2.664535259e-27   pdiblc1 = 0.39   pdiblc2 = 3.598389252e-04 lpdiblc2 = -5.862753804e-10   pdiblcb = -4.299292994e-04 lpdiblcb = -8.855717695e-9   drout = 0.56   pscbe1 = 7.804028631e+08 lpscbe1 = 7.932480083e+1   pscbe2 = 9.149943124e-09 lpscbe2 = 1.694800055e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -7.363294768e-01 lbeta0 = 3.006913896e-5   agidl = 1.924122583e-10 lagidl = -3.740640288e-16   bgidl = 7.993374236e+08 lbgidl = 1.614887265e+3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.109439203e-01 lkt1 = 4.458782848e-7   kt2 = -3.129229069e-02 lkt2 = -5.366827209e-8   at = -1.815528282e+05 lat = 1.461096312e+0   ute = 1.689857606e-01 lute = -4.013230319e-6   ua1 = 5.369873105e-09 lua1 = -2.310333602e-14   ub1 = -4.262076237e-18 lub1 = 2.077353037e-23   uc1 = 7.954823352e-10 luc1 = -2.974476434e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.043118709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.293769733e-7   k1 = 6.000718980e-01 lk1 = -3.259060697e-7   k2 = -9.796815934e-03 lk2 = 7.005882629e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.310204205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.376317553e-7   nfactor = {3.105619891e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.631739389e-6   eta0 = 0.08   etab = -0.07   u0 = 2.800388268e-03 lu0 = 1.353151645e-8   ua = -1.421659857e-09 lua = 1.962778754e-15   ub = 6.460886178e-19 lub = 1.180094484e-25   uc = -6.668216971e-11 luc = -3.764195286e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.460490681e+05 lvsat = -1.896466300e-1   a0 = 2.068078721e+00 la0 = -1.852248161e-6   ags = 5.238056873e-01 lags = -3.721365957e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -4.166157459e-02 lketa = 6.736539737e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.425310148e-01 lpclm = -1.253670861e-6   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = 2.029920012e-02 lpdiblcb = -9.276256952e-8   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.693071063e-08 lpscbe2 = -2.979999612e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.532589957e+00 lbeta0 = 4.693963595e-6   agidl = 1.0e-10   bgidl = 1.141376499e+09 lbgidl = 2.303900486e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.417866910e-01 lkt1 = -2.388321190e-7   kt2 = -4.004395473e-02 lkt2 = -1.824350515e-8   at = 2.774165791e+05 lat = -3.967085806e-1   ute = -1.664606991e+00 lute = 3.408740581e-6   ua1 = -3.361519923e-09 lua1 = 1.223937839e-14 pua1 = -1.323488980e-35   ub1 = 3.238276224e-18 lub1 = -9.586208816e-24 pub1 = 6.162975822e-45   uc1 = 9.309813477e-11 luc1 = -1.313832265e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.119082951e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.618070211e-8   k1 = 4.317830385e-01 lk1 = 1.871164947e-8   k2 = 2.813494163e-02 lk2 = -7.616878557e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 3.816385505e-01 ldsub = 3.652441172e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.107489027e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.563423735e-8   nfactor = {9.474016816e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.878059061e-7   eta0 = -6.563603097e-02 leta0 = 2.982298233e-7   etab = 7.292236481e-01 letab = -1.636630206e-06 petab = 1.332267630e-27   u0 = 1.047231551e-02 lu0 = -2.178864366e-9   ua = -1.340253773e-10 lua = -6.740069421e-16   ub = 4.537664404e-19 lub = 5.118419953e-25   uc = -1.236108384e-10 luc = 7.893515158e-17 wuc = -2.067951531e-31   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.960422668e+04 lvsat = 2.832845517e-2   a0 = 1.118388786e+00 la0 = 9.250314490e-8   ags = 9.605276213e-02 lags = 5.038051506e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -2.263989567e-03 lketa = -1.331199231e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.385327269e-02 lpclm = 6.275744520e-7   pdiblc1 = 4.099247304e-01 lpdiblc1 = -4.080136477e-8   pdiblc2 = -1.027162500e-05 lpdiblc2 = 4.613056019e-10   pdiblcb = -0.025   drout = 1.090551064e-01 ldrout = 9.234336795e-7   pscbe1 = 800000000.0   pscbe2 = -4.861149626e-09 lpscbe2 = 1.482483051e-14 ppscbe2 = -6.617444900e-36   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.732973460e+00 lbeta0 = 2.235848267e-6   agidl = 1.0e-10   bgidl = 1.269994274e+09 lbgidl = -3.299021648e+1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.436292395e-01 lkt1 = -3.028149435e-8   kt2 = -6.108811503e-02 lkt2 = 2.485020020e-08 wkt2 = 1.110223025e-22   at = 6.381357310e+04 lat = 4.070231495e-2   ute = 0.0   ua1 = 2.836786052e-09 lua1 = -4.533576282e-16   ub1 = -1.532069271e-18 lub1 = 1.823854303e-25   uc1 = 1.602296443e-10 luc1 = -2.688534535e-16 wuc1 = -1.033975766e-31 puc1 = -2.067951531e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.126492509e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.394425227e-8   k1 = 3.187815911e-01 lk1 = 1.371117410e-7   k2 = 6.539252981e-02 lk2 = -4.665444801e-08 wk2 = 5.551115123e-23   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 4.346808990e-01 ldsub = 3.096676706e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.878277982e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.618077084e-9   nfactor = {1.785445172e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.027511255e-8   eta0 = 3.750324212e-01 leta0 = -1.634915641e-7   etab = -1.744588252e+00 letab = 9.553680575e-7   u0 = 1.077941185e-02 lu0 = -2.500632234e-9   ua = -3.018047553e-10 lua = -4.982119042e-16   ub = 7.435590590e-19 lub = 2.082045343e-25   uc = -6.614406353e-11 luc = 1.872290159e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.907622725e+04 lvsat = 7.926179768e-3   a0 = 1.235349135e+00 la0 = -3.004498506e-8   ags = -1.637209281e-01 lags = 7.759895289e-7   a1 = 0.0   a2 = 5.809009555e-01 la2 = 2.295665014e-7   b0 = 0.0   b1 = 0.0   keta = 2.008093115e-02 lketa = -3.672444161e-08 pketa = -2.775557562e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.276496794e-01 lpclm = 9.970917197e-8   pdiblc1 = -3.181349608e-01 lpdiblc1 = 7.220413781e-7   pdiblc2 = -2.136988382e-04 lpdiblc2 = 6.744515502e-10   pdiblcb = -5.202309237e-02 lpdiblcb = 2.831412061e-8   drout = 1.011371724e+00 ldrout = -2.199111402e-8   pscbe1 = 8.095813297e+08 lpscbe1 = -1.003907775e+1   pscbe2 = 9.342690989e-09 lpscbe2 = -5.759858989e-17   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.412246329e+00 lbeta0 = 4.763481371e-7   agidl = 1.0e-10   bgidl = 1.285460944e+09 lbgidl = -4.919580623e+1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.518350605e-01 lkt1 = -2.168364023e-8   kt2 = -2.616352350e-02 lkt2 = -1.174291369e-8   at = 1.767849130e+05 lat = -7.766623072e-2   ute = 2.191100000e-02 lute = -2.295779803e-8   ua1 = 2.681055040e-09 lua1 = -2.901865670e-16   ub1 = -1.012244420e-18 lub1 = -3.622740528e-25   uc1 = -1.249950081e-10 luc1 = 2.999780679e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-9.689792327e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.233758270e-08 wvth0 = -1.639681155e-07 pvth0 = 8.981763447e-14   k1 = 2.163439841e+00 lk1 = -8.733459319e-07 wk1 = -3.332133355e-06 pk1 = 1.825259349e-12   k2 = -6.689544144e-01 lk2 = 3.556024493e-07 wk2 = 1.334571240e-06 pk2 = -7.310447611e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.350252821e+00 ldsub = -1.918597391e-07 wdsub = 2.765172429e-07 pdsub = -1.514692327e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.506992636e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.605749401e-08 wvoff = 1.880978919e-07 pvoff = -1.030353227e-13   nfactor = {2.066240048e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.440875255e-07 wnfactor = -1.869019096e-06 pnfactor = 1.023801935e-12   eta0 = -4.158717185e-01 leta0 = 2.697459510e-7   etab = -3.506512077e-04 letab = -8.169421162e-11   u0 = -3.696281518e-03 lu0 = 5.428790702e-09 wu0 = 1.938204162e-08 pu0 = -1.061699785e-14   ua = -3.961330771e-09 lua = 1.506384959e-15 wua = 5.780994451e-15 pua = -3.166684236e-21   ub = 2.334898557e-18 lub = -6.634914590e-25 wub = -3.264689430e-24 pub = 1.788315253e-30   uc = 2.061951598e-11 luc = -2.880401818e-17 wuc = -1.304958501e-16 puc = 7.148236427e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.604431599e+05 lvsat = -4.760009175e-02 wvsat = -1.838414392e-01 pvsat = 1.007037443e-7   a0 = 1.555335705e+00 la0 = -2.053256285e-07 wa0 = 2.073382178e-07 pa0 = -1.135746923e-13   ags = -6.039310850e+00 lags = 3.994490798e-06 wags = 1.179148735e-05 pags = -6.459081984e-12   a1 = 0.0   a2 = 4.132620724e-01 la2 = 3.213948905e-07 wa2 = 1.597267513e-06 pa2 = -8.749432121e-13   b0 = 0.0   b1 = 0.0   keta = -5.750673288e-02 lketa = 5.776141051e-09 wketa = 6.726843540e-08 pketa = -3.684796720e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.372507777e+00 lpclm = -3.630829727e-07 wpclm = -1.119446950e-06 ppclm = 6.132050532e-13   pdiblc1 = 2.248484686e+00 lpdiblc1 = -6.838886987e-07 wpdiblc1 = -9.812480307e-07 ppdiblc1 = 5.375031400e-13   pdiblc2 = 3.888965943e-03 lpdiblc2 = -1.572885650e-09 wpdiblc2 = -2.170076990e-08 ppdiblc2 = 1.188713923e-14   pdiblcb = -1.171829384e+00 lpdiblcb = 6.417160121e-07 wpdiblcb = 2.325173704e-06 ppdiblcb = -1.273672026e-12   drout = 3.085850619e+00 ldrout = -1.158338791e-06 wdrout = -2.865584856e-06 pdrout = 1.569695745e-12   pscbe1 = 7.818992258e+08 lpscbe1 = 5.124486733e+00 wpscbe1 = -1.716253895e+00 ppscbe1 = 9.401209772e-7   pscbe2 = 1.043059010e-08 lpscbe2 = -6.535225257e-16 wpscbe2 = -2.086950477e-15 ppscbe2 = 1.143179297e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.133553993e+01 lbeta0 = -1.124959014e-06 wbeta0 = -2.673449986e-06 pbeta0 = 1.464449066e-12   agidl = 1.426811023e-09 lagidl = -7.267939079e-16 wagidl = -2.569013960e-15 pagidl = 1.407241622e-21   bgidl = 1.141474556e+09 lbgidl = 2.967633718e+01 wbgidl = 4.642072406e+02 pbgidl = -2.542811212e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -6.564357404e-01 lkt1 = 9.039149719e-08 wkt1 = 3.137915042e-07 pkt1 = -1.718871412e-13   kt2 = -3.816507159e-02 lkt2 = -5.168765683e-09 wkt2 = -1.295786354e-08 pkt2 = 7.097993700e-15   at = -1.801252157e+05 lat = 1.178402150e-01 wat = 3.960691057e-01 pat = -2.169567544e-7   ute = -1.641403659e-01 lute = 7.895648895e-08 wute = 2.329642703e-07 pute = -1.276120032e-13   ua1 = -2.983016966e-09 lua1 = 2.812450476e-15 wua1 = 1.079686519e-14 pua1 = -5.914252830e-21   ub1 = 3.917236481e-18 lub1 = -3.062520453e-24 wub1 = -1.135476812e-23 pub1 = 6.219858108e-30   uc1 = 5.340306734e-10 luc1 = -3.309999859e-16 wuc1 = -1.061276983e-15 puc1 = 5.813409994e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.421891802e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.252845752e-08 wvth0 = 5.856004125e-07 pvth0 = -1.333851340e-13   k1 = -6.401670772e+00 lk1 = 1.677129881e-06 wk1 = 1.190047627e-05 pk1 = -2.710630982e-12   k2 = 2.781029817e+00 lk2 = -6.717166052e-07 wk2 = -4.766325858e-06 pk2 = 1.085649872e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.173330524e+00 ldsub = -1.391767019e-07 wdsub = -9.875615819e-07 pdsub = 2.249418393e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {1.883266935e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.467346035e-08 wvoff = -6.717781853e-07 pvoff = 1.530142762e-13   nfactor = {-1.912611464e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.407149834e-07 wnfactor = 6.675068199e-06 pnfactor = -1.520413659e-12   eta0 = 0.49   etab = -0.000625   u0 = 4.729578605e-02 lu0 = -9.755372218e-09 wu0 = -6.922157722e-08 pu0 = 1.576694475e-14   ua = 1.086891351e-08 lua = -2.909691031e-15 wua = -2.064640875e-14 pua = 4.702735754e-21   ub = -5.411471869e-18 lub = 1.643183994e-24 wub = 1.165960511e-23 pub = -2.655766554e-30   uc = -2.966845217e-10 luc = 6.568119165e-17 wuc = 4.660566074e-16 puc = -1.061560437e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -3.101510594e+05 lvsat = 9.253110190e-02 wvsat = 6.565765685e-01 pvsat = -1.495517279e-7   a0 = 1.216260483e+00 la0 = -1.043575042e-07 wa0 = -7.404936351e-07 pa0 = 1.686659377e-13   ags = 2.730594666e+01 lags = -5.934893257e-06 wags = -4.211245483e-05 pags = 9.592164398e-12   a1 = 0.0   a2 = 4.192396738e+00 la2 = -8.039369345e-07 wa2 = -5.704526833e-06 pa2 = 1.299348599e-12   b0 = 0.0   b1 = 0.0   keta = 7.559275657e-02 lketa = -3.385755942e-08 wketa = -2.402444121e-07 pketa = 5.472167097e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.738979710e+00 lpclm = 5.634402140e-07 wpclm = 3.998024823e-06 ppclm = -9.106501040e-13   pdiblc1 = -1.706752023e+00 lpdiblc1 = 4.938819122e-07 wpdiblc1 = 3.504457252e-06 ppdiblc1 = -7.982277507e-13   pdiblc2 = -3.807332285e-02 lpdiblc2 = 1.092243490e-08 wpdiblc2 = 7.750274963e-08 ppdiblc2 = -1.765318880e-14   pdiblcb = 4.913378590e+00 lpdiblcb = -1.170306792e-06 wpdiblcb = -8.304191802e-06 ppdiblcb = 1.891487288e-12   drout = -5.647741552e+00 ldrout = 1.442306618e-06 wdrout = 1.023423163e-05 pdrout = -2.331102109e-12   pscbe1 = 7.962075510e+08 lpscbe1 = 8.638251786e-01 wpscbe1 = 6.129478196e+00 ppscbe1 = -1.396141896e-6   pscbe2 = 4.708394598e-09 lpscbe2 = 1.050404240e-15 wpscbe2 = 7.453394560e-15 ppscbe2 = -1.697696946e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.038804880e+00 lbeta0 = 1.345601265e-06 wbeta0 = 9.548035663e-06 pbeta0 = -2.174803823e-12   agidl = -5.356264843e-09 lagidl = 1.293036508e-15 wagidl = 9.175049857e-15 pagidl = -2.089846981e-21   bgidl = 2.025770411e+09 lbgidl = -2.336448609e+02 wbgidl = -1.657883002e+03 pbgidl = 3.776243008e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 1.775129999e-01 lkt1 = -1.579375889e-07 wkt1 = -1.120683944e-06 pkt1 = 2.552637852e-13   kt2 = -7.742531703e-02 lkt2 = 6.521953902e-09 wkt2 = 4.627808407e-08 pkt2 = -1.054099060e-14   at = 8.850742779e+05 lat = -1.993495642e-01 wat = -1.414532520e+00 pat = 3.221951448e-7   ute = 4.947870185e-01 lute = -1.172556129e-07 wute = -8.320152511e-07 pute = 1.895122738e-13   ua1 = 2.471148510e-08 lua1 = -5.434279875e-15 wua1 = -3.856023282e-14 pua1 = 8.783057031e-21   ub1 = -2.556006725e-17 lub1 = 5.715083666e-24 wub1 = 4.055274329e-23 pub1 = -9.236901104e-30   uc1 = -2.371391484e-09 luc1 = 5.341620970e-16 wuc1 = 3.790274940e-15 puc1 = -8.633298744e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.169233938e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.684364501e-08 wvth0 = 2.129737799e-07 pvth0 = -5.213065699e-14   k1 = 1.897196960e-01 lk1 = 1.888949626e-07 wk1 = -2.267541197e-07 pk1 = 5.550373965e-14   k2 = 1.492419512e-01 lk2 = -7.765433710e-08 wk2 = 5.546035477e-08 pk2 = -1.357530834e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.645676761e+00 ldsub = -5.099577131e-07 wdsub = -2.843889120e-07 pdsub = 6.961129595e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {2.119901634e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.083074225e-08 wvoff = -5.018037322e-07 pvoff = 1.228290085e-13   nfactor = {1.682484377e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.575535305e-06 wnfactor = -2.325832664e-05 pnfactor = 5.693056904e-12   eta0 = -2.673913572e-02 leta0 = 1.264848219e-07 weta0 = 4.743473667e-06 peta0 = -1.161083767e-12   etab = -1.628074271e+00 letab = 3.983588953e-07 wetab = 3.148603298e-06 petab = -7.706993723e-13   u0 = 3.407008347e-02 lu0 = -7.246143625e-09 wu0 = -4.777981546e-08 pu0 = 1.169530433e-14   ua = 1.297299343e-08 lua = -3.641882149e-15 wua = -2.563852363e-14 pua = 6.275669621e-21   ub = -1.257474851e-17 lub = 3.519214164e-24 wub = 2.580942250e-23 pub = -6.317501392e-30   uc = -7.094416139e-11 luc = 1.532771440e-17 wuc = 1.417892877e-16 puc = -3.470647290e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.535390646e+05 lvsat = -1.119725842e-01 wvsat = -3.011233199e-01 pvsat = 7.370746063e-8   a0 = -9.188376287e+00 la0 = 2.434648733e-06 wa0 = 1.728670524e-05 pa0 = -4.231353276e-12   ags = 1.249999777e+00 lags = 4.780483565e-14   a1 = 0.0   a2 = -2.295741368e+00 la2 = 7.241951919e-07 wa2 = 4.367621014e-06 pa2 = -1.069084434e-12   b0 = 7.619782290e-23 lb0 = -1.865132210e-29 wb0 = -1.475366630e-28 pb0 = 3.611328669e-35   b1 = 0.0   keta = -7.770173487e-01 lketa = 1.723131182e-07 wketa = 4.978556938e-07 pketa = -1.218626275e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.866249091e+00 lpclm = -5.217522736e-07 wpclm = -2.657124199e-06 ppclm = 6.503975757e-13   pdiblc1 = 2.828728472e+00 lpdiblc1 = -5.794294215e-07 wpdiblc1 = -4.071879537e-07 ppdiblc1 = 9.966943138e-14   pdiblc2 = 7.384293986e-02 lpdiblc2 = -1.565667176e-08 wpdiblc2 = -3.545590563e-08 ppdiblc2 = 8.678719301e-15   pdiblcb = 4.479745766e+01 lpdiblcb = -1.102027816e-05 wpdiblcb = -7.449730840e-05 ppdiblcb = 1.823507866e-11   drout = -1.574920319e+00 ldrout = 5.530284364e-07 wdrout = -4.045213416e-12 pdrout = 9.901671127e-19   pscbe1 = 7.864931781e+08 lpscbe1 = 3.306132464e+00 wpscbe1 = 2.615234903e+01 ppscbe1 = -6.401441234e-6   pscbe2 = -4.604878288e-08 lpscbe2 = 1.355288934e-14 wpscbe2 = 1.074823457e-13 ppscbe2 = -2.630899117e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 2.323404954e+01 lbeta0 = -3.497260719e-06 wbeta0 = -1.509249330e-05 pbeta0 = 3.694265048e-12   agidl = 2.118532789e-08 lagidl = -5.107176000e-15 wagidl = -3.777172009e-14 pagidl = 9.245572786e-21   bgidl = 9.999997992e+08 lbgidl = 4.312079430e-5   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.717525279e-01 lkt1 = 1.367619975e-08 wkt1 = 4.200729771e-07 pkt1 = -1.028233630e-13   kt2 = -1.765666763e-02 lkt2 = -7.621150857e-09 wkt2 = -1.816818194e-13 pkt2 = 4.447116742e-20   at = 2.257898459e+05 lat = -5.285168332e-02 wat = -5.734000178e-01 pat = 1.403539894e-7   ute = 1.834223514e+00 lute = -4.538675605e-07 wute = 1.065690369e-12 pute = -2.608543607e-19   ua1 = 6.140093501e-09 lua1 = -1.294055283e-15 wua1 = -4.200732891e-15 pua1 = 1.028234393e-21   ub1 = -2.813062721e-18 lub1 = 5.737312242e-25 wub1 = 1.859445807e-30 pub1 = -4.551458486e-37   uc1 = -9.741274361e-10 luc1 = 2.320140080e-16 wuc1 = 1.834319069e-15 puc1 = -4.489954501e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.094269313e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.397621949e-8   k1 = 4.212225495e-01 lk1 = 1.296244034e-06 wk1 = -7.105427358e-21   k2 = 4.426361306e-02 lk2 = -5.789263560e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.795342868e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.623402023e-7   nfactor = {1.120644890e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.684324920e-5   eta0 = 0.08   etab = -0.07   u0 = 9.292746448e-03 lu0 = -1.593665493e-8   ua = -6.110105453e-11 lua = -4.383983995e-15 pua = -2.646977960e-35   ub = 7.489433296e-20 lub = 3.936931675e-24   uc = -7.212777231e-11 luc = -7.432635937e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160312.5   a0 = 1.750746838e+00 la0 = -2.073473977e-6   ags = 4.164861845e-01 lags = 3.191979779e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -5.481686414e-02 lketa = 4.727443598e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.043571226e-01 lpclm = -2.891108831e-6   pdiblc1 = 0.39   pdiblc2 = 1.361647904e-04 lpdiblc2 = 3.023700845e-9   pdiblcb = -3.449935132e-03 lpdiblcb = 3.848396013e-8   drout = 0.56   pscbe1 = 7.008212287e+08 lpscbe1 = 1.793040344e+3   pscbe2 = 9.666159942e-09 lpscbe2 = -6.127090055e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 5.684079876e-10 lalpha0 = -9.390537943e-15   alpha1 = -2.471546770e-11 lalpha1 = 2.500267635e-15 walpha1 = -3.877409121e-32 palpha1 = 1.344168495e-36   beta0 = 3.268606140e+00 lbeta0 = -5.384955464e-6   agidl = 8.848961259e-11 lagidl = 1.151588650e-15   bgidl = 1.563280604e+09 lbgidl = -1.129252281e+4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.257132571e-01 lkt1 = -5.979598311e-7   kt2 = -0.037961   at = 0.0   ute = -3.560025648e-01 lute = 5.275083793e-7   ua1 = 2.139553309e-09 lua1 = 7.208111171e-15   ub1 = -7.300459942e-19 lub1 = -1.906050239e-23   uc1 = 4.315974271e-11 luc1 = 7.672689606e-15 puc1 = -5.293955920e-35   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.0895817+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.4858803   k2 = 0.015386276   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.17143662+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.4596089+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.0084978126   ua = -2.7977789e-10   ub = 2.7127182e-19   uc = -1.0920239e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160312.5   a0 = 1.6473202   ags = 0.43240805   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -0.031235975   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.060146165   pdiblc1 = 0.39   pdiblc2 = 0.00028698955   pdiblcb = -0.0015303226   drout = 0.56   pscbe1 = 790259600.0   pscbe2 = 9.3605355e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.0   agidl = 1.4593183e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.45554   kt2 = -0.037961   at = 0.0   ute = -0.32969   ua1 = 2.4991e-9   ub1 = -1.6808e-18   uc1 = 4.2588e-10   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.104255390e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.180905583e-7   k1 = 4.518013436e-01 lk1 = 2.742597737e-7   k2 = 2.335544192e-02 lk2 = -6.413405423e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.779276016e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.223795970e-8   nfactor = {2.713816962e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.045809286e-6   eta0 = 0.08   etab = -0.07   u0 = 1.088040643e-02 lu0 = -1.917457908e-8   ua = 3.850477410e-10 lua = -5.350367093e-15   ub = -1.375240580e-19 lub = 3.289897247e-24   uc = -1.428199730e-10 luc = 2.705467437e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.221579483e+05 lvsat = -4.977182523e-1   a0 = 1.684598285e+00 la0 = -3.000056410e-7   ags = 4.329529311e-01 lags = -4.385080593e-9   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -3.752720400e-02 lketa = 5.063039543e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.193599535e-01 lpclm = 4.663734853e-06 wpclm = -1.776356839e-21 ppclm = -1.421085472e-26   pdiblc1 = 0.39   pdiblc2 = 3.598389252e-04 lpdiblc2 = -5.862753804e-10   pdiblcb = -4.299292994e-04 lpdiblcb = -8.855717695e-9   drout = 0.56   pscbe1 = 7.804028631e+08 lpscbe1 = 7.932480083e+1   pscbe2 = 9.149943124e-09 lpscbe2 = 1.694800055e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -7.363294768e-01 lbeta0 = 3.006913896e-5   agidl = 1.924122583e-10 lagidl = -3.740640288e-16   bgidl = 7.993374236e+08 lbgidl = 1.614887265e+3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.109439203e-01 lkt1 = 4.458782848e-7   kt2 = -3.129229069e-02 lkt2 = -5.366827209e-8   at = -1.815528282e+05 lat = 1.461096312e+0   ute = 1.689857606e-01 lute = -4.013230319e-6   ua1 = 5.369873105e-09 lua1 = -2.310333602e-14 pua1 = 2.117582368e-34   ub1 = -4.262076237e-18 lub1 = 2.077353037e-23 wub1 = -4.930380658e-38   uc1 = 7.954823353e-10 luc1 = -2.974476434e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.043118709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.293769733e-7   k1 = 6.000718980e-01 lk1 = -3.259060697e-7   k2 = -9.796815934e-03 lk2 = 7.005882629e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.310204205e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.376317553e-7   nfactor = {3.105619891e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.631739389e-6   eta0 = 0.08   etab = -0.07   u0 = 2.800388268e-03 lu0 = 1.353151645e-8   ua = -1.421659857e-09 lua = 1.962778754e-15   ub = 6.460886178e-19 lub = 1.180094484e-25   uc = -6.668216971e-11 luc = -3.764195286e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.460490681e+05 lvsat = -1.896466300e-1   a0 = 2.068078721e+00 la0 = -1.852248161e-6   ags = 5.238056873e-01 lags = -3.721365957e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -4.166157459e-02 lketa = 6.736539737e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.425310148e-01 lpclm = -1.253670861e-6   pdiblc1 = 0.39   pdiblc2 = 0.000215   pdiblcb = 2.029920012e-02 lpdiblcb = -9.276256952e-08 wpdiblcb = -5.551115123e-23   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.693071063e-08 lpscbe2 = -2.979999612e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.532589957e+00 lbeta0 = 4.693963595e-6   agidl = 1.0e-10   bgidl = 1.141376499e+09 lbgidl = 2.303900486e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.417866910e-01 lkt1 = -2.388321190e-7   kt2 = -4.004395473e-02 lkt2 = -1.824350515e-8   at = 2.774165791e+05 lat = -3.967085806e-1   ute = -1.664606991e+00 lute = 3.408740581e-6   ua1 = -3.361519923e-09 lua1 = 1.223937839e-14 wua1 = 1.323488980e-29 pua1 = 1.058791184e-34   ub1 = 3.238276224e-18 lub1 = -9.586208816e-24 pub1 = 4.930380658e-44   uc1 = 9.309813477e-11 luc1 = -1.313832265e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.119082951e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.618070211e-8   k1 = 4.317830385e-01 lk1 = 1.871164947e-8   k2 = 2.813494163e-02 lk2 = -7.616878557e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 3.816385505e-01 ldsub = 3.652441172e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.107489027e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.563423735e-8   nfactor = {9.474016816e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.878059061e-7   eta0 = -6.563603097e-02 leta0 = 2.982298233e-7   etab = 7.292236481e-01 letab = -1.636630206e-06 wetab = -3.552713679e-21 petab = -1.065814104e-26   u0 = 1.047231551e-02 lu0 = -2.178864366e-9   ua = -1.340253773e-10 lua = -6.740069421e-16   ub = 4.537664404e-19 lub = 5.118419953e-25   uc = -1.236108384e-10 luc = 7.893515158e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.960422668e+04 lvsat = 2.832845517e-2   a0 = 1.118388786e+00 la0 = 9.250314490e-8   ags = 9.605276213e-02 lags = 5.038051506e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -2.263989567e-03 lketa = -1.331199231e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.385327269e-02 lpclm = 6.275744520e-7   pdiblc1 = 4.099247304e-01 lpdiblc1 = -4.080136477e-8   pdiblc2 = -1.027162500e-05 lpdiblc2 = 4.613056019e-10   pdiblcb = -0.025   drout = 1.090551064e-01 ldrout = 9.234336795e-7   pscbe1 = 800000000.0   pscbe2 = -4.861149626e-09 lpscbe2 = 1.482483051e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.732973460e+00 lbeta0 = 2.235848267e-6   agidl = 1.0e-10   bgidl = 1.269994274e+09 lbgidl = -3.299021648e+1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.436292395e-01 lkt1 = -3.028149435e-8   kt2 = -6.108811503e-02 lkt2 = 2.485020020e-8   at = 6.381357310e+04 lat = 4.070231495e-2   ute = 0.0   ua1 = 2.836786052e-09 lua1 = -4.533576282e-16   ub1 = -1.532069271e-18 lub1 = 1.823854303e-25   uc1 = 1.602296443e-10 luc1 = -2.688534535e-16 wuc1 = 8.271806126e-31 puc1 = -8.271806126e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.126492509e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.394425227e-8   k1 = 3.187815911e-01 lk1 = 1.371117410e-7   k2 = 6.539252981e-02 lk2 = -4.665444801e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 4.346808990e-01 ldsub = 3.096676706e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.878277982e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.618077084e-9   nfactor = {1.785445172e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.027511255e-8   eta0 = 3.750324212e-01 leta0 = -1.634915641e-07 weta0 = -7.105427358e-21   etab = -1.744588252e+00 letab = 9.553680575e-7   u0 = 1.077941185e-02 lu0 = -2.500632234e-9   ua = -3.018047553e-10 lua = -4.982119042e-16   ub = 7.435590590e-19 lub = 2.082045343e-25   uc = -6.614406353e-11 luc = 1.872290159e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.907622725e+04 lvsat = 7.926179768e-3   a0 = 1.235349135e+00 la0 = -3.004498506e-8   ags = -1.637209281e-01 lags = 7.759895289e-7   a1 = 0.0   a2 = 5.809009555e-01 la2 = 2.295665014e-7   b0 = 0.0   b1 = 0.0   keta = 2.008093115e-02 lketa = -3.672444161e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.276496794e-01 lpclm = 9.970917197e-8   pdiblc1 = -3.181349608e-01 lpdiblc1 = 7.220413781e-7   pdiblc2 = -2.136988382e-04 lpdiblc2 = 6.744515502e-10   pdiblcb = -5.202309237e-02 lpdiblcb = 2.831412061e-8   drout = 1.011371724e+00 ldrout = -2.199111402e-8   pscbe1 = 8.095813297e+08 lpscbe1 = -1.003907775e+1   pscbe2 = 9.342690989e-09 lpscbe2 = -5.759858989e-17   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.412246329e+00 lbeta0 = 4.763481371e-7   agidl = 1.0e-10   bgidl = 1.285460944e+09 lbgidl = -4.919580623e+1   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.518350605e-01 lkt1 = -2.168364023e-8   kt2 = -2.616352350e-02 lkt2 = -1.174291369e-8   at = 1.767849130e+05 lat = -7.766623072e-2   ute = 2.191100000e-02 lute = -2.295779803e-8   ua1 = 2.681055040e-09 lua1 = -2.901865670e-16   ub1 = -1.012244420e-18 lub1 = -3.622740528e-25   uc1 = -1.249950081e-10 luc1 = 2.999780679e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.070430086e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.234658453e-9   k1 = 1.017721134e-01 lk1 = 2.559841077e-7   k2 = 1.567755799e-01 lk2 = -9.671179828e-08 wk2 = 4.440892099e-22 pk2 = 2.220446049e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.521340414e+00 ldsub = -2.855772454e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.343187613e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.769283561e-8   nfactor = {9.098348438e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.893623352e-7   eta0 = -4.158717185e-01 leta0 = 2.697459510e-07 weta0 = -3.552713679e-21 peta0 = -8.881784197e-28   etab = -3.506512077e-04 letab = -8.169421162e-11   u0 = 8.295834478e-03 lu0 = -1.140190638e-9   ua = -3.844962256e-10 lua = -4.529155841e-16   ub = 3.149599400e-19 lub = 4.429804168e-25   uc = -6.012127499e-11 luc = 1.542376859e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 4.669622306e+04 lvsat = 1.470763656e-2   a0 = 1.683620641e+00 la0 = -2.755969091e-7   ags = 1.256354222e+00 lags = -1.892136726e-9   a1 = 0.0   a2 = 1.401528307e+00 la2 = -2.199526463e-7   b0 = 0.0   b1 = 0.0   keta = -1.588620105e-02 lketa = -1.702254577e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.798801408e-01 lpclm = 1.632113096e-8   pdiblc1 = 1.641363907e+00 lpdiblc1 = -3.513231140e-7   pdiblc2 = -9.537800695e-03 lpdiblc2 = 5.781961445e-09 wpdiblc2 = -2.775557562e-23 ppdiblc2 = 2.081668171e-29   pdiblcb = 2.668091928e-01 lpdiblcb = -1.463342344e-07 wpdiblcb = 8.118505868e-22 ppdiblcb = -6.661338148e-28   drout = 1.312847203e+00 ldrout = -1.871318449e-7   pscbe1 = 7.808373399e+08 lpscbe1 = 5.706161256e+0   pscbe2 = 9.139345727e-09 lpscbe2 = 5.378886116e-17   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.681414786e+00 lbeta0 = -2.188706146e-7   agidl = -1.626971420e-10 lagidl = 1.438989270e-16 pagidl = 8.271806126e-37   bgidl = 1.428690278e+09 lbgidl = -1.276532549e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.622857024e-01 lkt1 = -1.595903986e-8   kt2 = -4.618240050e-02 lkt2 = -7.770733397e-10   at = 6.493187118e+04 lat = -1.639593073e-2   ute = -2.000000099e-02 lute = 5.447382545e-16   ua1 = 3.697252445e-09 lua1 = -8.468341008e-16   ub1 = -3.108220336e-18 lub1 = 7.858491546e-25 pub1 = -1.232595164e-44   uc1 = -1.226058634e-10 luc1 = 2.868909302e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.05956732562893+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.961428255393082   k2 = -0.168005876831761   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.562303405039308   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.227317957389937+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.2174071222327+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.49   etab = -0.000625   u0 = 0.0044668003490566   ua = -1.90549558459119e-9   ub = 1.80259461966667e-18   uc = -8.324553995283e-12   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 96088.000620792   a0 = 0.758099999261006   ags = 1.24999997272013   a1 = 0.0   a2 = 0.662874470440252   b0 = 0.0   b1 = 0.0   keta = -0.0730519999606918   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.734690420259434   pdiblc1 = 0.461536473183962   pdiblc2 = 0.00987941513820755   pdiblcb = -0.224616327814465   drout = 0.684413503600629   pscbe1 = 800000000.518868   pscbe2 = 9.31998164677673e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.94639467130503   agidl = 3.20550031084906e-10   bgidl = 999999975.393082   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.515879992940252   kt2 = -0.0487919994941038   at = 9870.39612421382   ute = -0.0199999991650943   ua1 = 8.53380055896226e-10   ub1 = -4.69150049528303e-19   uc1 = -2.62609955581761e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.037445128e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.414960836e-09 wvth0 = -2.751122838e-11 pvth0 = 6.734060946e-18   k1 = 4.942515946e-02 lk1 = 2.232355578e-07 wk1 = -5.600377790e-12 pk1 = 1.370832479e-18   k2 = 1.835509467e-01 lk2 = -8.605232149e-08 wk2 = 9.058230319e-12 pk2 = -2.217228321e-18   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.469696404e+00 ldsub = -4.668821214e-07 wdsub = 3.617126498e-11 pdsub = -8.853821370e-18   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.892779319e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.516625277e-08 wvoff = -9.530924672e-13 pvoff = 2.332932070e-19   nfactor = {2.434364820e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.310582037e-08 wnfactor = 2.592744772e-11 pnfactor = -6.346390990e-18   eta0 = 2.908147341e+00 leta0 = -5.919020153e-07 weta0 = 1.622697363e-11 peta0 = -3.971957469e-18   etab = 3.200414198e-01 letab = -7.849112290e-08 wetab = -3.620851520e-12 petab = 8.862939306e-19   u0 = 4.507584642e-03 lu0 = -9.982975393e-12 wu0 = 4.114224250e-14 pu0 = -1.007059247e-20   ua = -2.890138196e-09 lua = 2.410158952e-16 wua = -2.267126691e-20 pua = 5.549359330e-27   ub = 3.394140339e-18 lub = -3.895706034e-25 wub = -6.663942334e-30 pub = 1.631166447e-36   uc = 1.678410277e-11 luc = -6.145971460e-18 wuc = 5.985727977e-23 puc = -1.465156564e-29   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.672317794e+05 lvsat = -6.636921845e-02 wvsat = -7.523805104e-06 pvsat = 1.841639396e-12   a0 = 1.507303731e+00 la0 = -1.833863433e-07 wa0 = 4.937583299e-12 pa0 = -1.208596956e-18   ags = 1.249999777e+00 lags = 4.780483209e-14   a1 = 0.0   a2 = 4.065942930e-01 la2 = 6.273098043e-08 wa2 = 1.964371984e-11 pa2 = -4.808291521e-18   b0 = -1.508642251e-23 lb0 = 3.692779069e-30 wb0 = -1.445052274e-34 pb0 = 3.537126707e-41   b1 = 0.0   keta = -4.689806504e-01 lketa = 9.691343541e-08 wketa = -3.075071326e-12 pketa = 7.527005845e-19   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.222227336e+00 lpclm = -1.193368485e-07 wpclm = -3.629072353e-12 ppclm = 8.883062037e-19   pdiblc1 = 2.576802988e+00 lpdiblc1 = -5.177643612e-07 wpdiblc1 = -1.792507089e-11 ppdiblc1 = 4.387609209e-18   pdiblc2 = 5.190541848e-02 lpdiblc2 = -1.028691497e-08 wpdiblc2 = 2.184276813e-13 ppdiblc2 = -5.346563570e-20   pdiblcb = -1.295745055e+00 lpdiblcb = 2.621855343e-07 wpdiblcb = 8.092293626e-13 ppdiblcb = -1.980791211e-19   drout = -1.574944693e+00 ldrout = 5.530344026e-07 wdrout = 3.534919074e-11 pdrout = -8.652598154e-18   pscbe1 = 8.026732801e+08 lpscbe1 = -6.543520080e-01 wpscbe1 = 1.550380493e-03 ppscbe1 = -3.794943848e-10   pscbe2 = 2.045293512e-08 lpscbe2 = -2.725068687e-15 wpscbe2 = 1.410114108e-19 ppscbe2 = -3.451606786e-26   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.389599333e+01 lbeta0 = -1.211538013e-06 wbeta0 = -2.805071017e-11 pbeta0 = 6.866112699e-18   agidl = -2.184899364e-09 lagidl = 6.132713757e-16 wagidl = -1.096569939e-20 pagidl = 2.684129077e-27   bgidl = 9.999997992e+08 lbgidl = 4.312080383e-5   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.118429970e-01 lkt1 = -4.994315568e-08 wkt1 = -1.123929849e-12 pkt1 = 2.751099402e-19   kt2 = -1.765776234e-02 lkt2 = -7.620882899e-09 wkt2 = 1.587630770e-12 pkt2 = -3.886123219e-19   at = -1.289843648e+05 lat = 3.398817411e-02 wat = -2.585680231e-06 pat = 6.329098779e-13   ute = 1.834229935e+00 lute = -4.538691322e-07 wute = -9.312559881e-12 pute = 2.279481840e-18   ua1 = 3.540999257e-09 lua1 = -6.578619898e-16 wua1 = 6.396764760e-21 pua1 = -1.565768090e-27   ub1 = -2.813051517e-18 lub1 = 5.737284818e-25 wub1 = -1.624881010e-29 pub1 = 3.977302491e-36   uc1 = 1.608061745e-10 luc1 = -4.578936656e-17 wuc1 = 3.049381476e-21 puc1 = -7.464123500e-28   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.128142877e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.332699994e-06 wvth0 = 5.373133081e-08 pvth0 = -3.551135290e-12   k1 = 1.934130088e-01 lk1 = 8.222303209e-06 wk1 = 3.613587834e-07 pk1 = -1.098633670e-11   k2 = 1.356026544e-01 lk2 = -2.631246592e-06 wk2 = -1.448849103e-07 pk2 = 3.255456033e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.288251500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.106768439e-06 wvoff = 7.818674456e-08 pvoff = -4.670546290e-12   nfactor = {-3.519184828e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.624916643e-04 wnfactor = 7.359846374e-06 pnfactor = -2.151698568e-10   eta0 = 0.08   etab = -0.07   u0 = 1.300734532e-02 lu0 = -1.925124052e-07 wu0 = -5.892215591e-09 pu0 = 2.800901055e-13   ua = 2.803433038e-10 lua = 1.511439141e-14 wua = -5.416099674e-16 pua = -3.092894702e-20   ub = 2.773646358e-19 lub = -6.450706067e-23 wub = -3.211648734e-25 pub = 1.085680509e-28   uc = 7.035676458e-11 luc = -5.901120570e-15 wuc = -2.260135319e-16 puc = 8.181557787e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.603105784e+05 lvsat = 1.922535840e-04 wvsat = 3.048131626e-06 pvsat = -3.049587871e-10   a0 = 1.734512602e+00 la0 = 2.492964928e-05 wa0 = 2.575126531e-08 pa0 = -4.283321821e-11   ags = 2.518921334e-01 lags = 1.287954450e-05 wags = 2.610843508e-07 pags = -1.992362359e-11   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -1.045737002e-01 lketa = -3.354952443e-07 wketa = 7.892588560e-08 pketa = 1.282055524e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 7.088063835e-01 lpclm = -1.797351708e-05 wpclm = -8.001735600e-07 ppclm = 2.392419860e-11   pdiblc1 = 0.39   pdiblc2 = -3.016203816e-04 lpdiblc2 = 9.813614491e-09 wpdiblc2 = 6.944288489e-10 ppdiblc2 = -1.077037830e-14   pdiblcb = -1.273937900e-01 lpdiblcb = 1.196775457e-05 wpdiblcb = 1.966037087e-07 ppdiblcb = -1.892259077e-11   drout = 0.56   pscbe1 = 4.339398113e+08 lpscbe1 = 6.547462248e+03 wpscbe1 = 4.233358446e+02 ppscbe1 = -7.541616166e-3   pscbe2 = 7.578907762e-09 lpscbe2 = 2.776922542e-13 wpscbe2 = 3.310866201e-15 ppscbe2 = -4.502033261e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.005137792e-09 lalpha0 = -3.819377380e-14 walpha0 = -2.278986791e-15 palpha0 = 4.568861442e-20   alpha1 = -4.072504250e-10 lalpha1 = 1.016924239e-14 walpha1 = 6.067891904e-16 palpha1 = -1.216477316e-20   beta0 = 6.612569630e+00 lbeta0 = -2.740302396e-04 wbeta0 = -5.304301894e-06 pbeta0 = 4.261337464e-10   agidl = 1.422523143e-10 lagidl = -1.832247437e-14 wagidl = -8.528011791e-17 pagidl = 3.089038193e-20   bgidl = 3.291009535e+09 lbgidl = -4.592964368e+04 wbgidl = -2.740578918e+03 pbgidl = 5.494250952e-2   cgidl = 300.0   egidl = 7.037336073e-01 legidl = -6.040220411e-05 wegidl = -9.576615674e-07 pegidl = 9.581190903e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.228750708e-01 lkt1 = -3.567777845e-06 wkt1 = -1.631252219e-07 pkt1 = 4.710820367e-12   kt2 = -4.902757531e-02 lkt2 = 1.107186237e-06 wkt2 = 1.755415589e-08 pkt2 = -1.756254239e-12   at = 0.0   ute = -2.849607871e-01 lute = -1.303666486e-05 wute = -1.126887411e-07 pute = 2.151592564e-11   ua1 = 5.168353404e-10 lua1 = 8.133153432e-14 wua1 = 2.574007168e-15 pua1 = -1.175769457e-19   ub1 = 2.927841349e-18 lub1 = -1.517270967e-22 wub1 = -5.802257956e-24 pub1 = 2.104399972e-28   uc1 = -1.464829142e-09 luc1 = 6.463137223e-14 wuc1 = 2.392020225e-15 puc1 = -9.034968505e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.011785825e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.234023057e-7   k1 = 6.035484582e-01 wk1 = -1.866489979e-7   k2 = 4.353845412e-03 wk2 = 1.749999444e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-7.385690850e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = -1.547840609e-7   nfactor = {4.586037038e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -3.373008358e-6   eta0 = 0.08   etab = -0.07   u0 = 3.404663463e-03 wu0 = 8.078916142e-9   ua = 1.034261951e-09 wua = -2.084372045e-15   ub = -2.940302196e-18 wub = 5.094301475e-24   uc = -2.239961284e-10 wuc = 1.820895013e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.603201682e+05 wvsat = -1.216347101e-5   a0 = 2.978024627e+00 wa0 = -2.110805944e-6   ags = 8.943347238e-01 wags = -7.327228716e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -1.213084872e-01 wketa = 1.428759012e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.877278743e-01 wpclm = 3.931857331e-7   pdiblc1 = 0.39   pdiblc2 = 1.878910226e-04 wpdiblc2 = 1.571932553e-10   pdiblcb = 4.695679460e-01 wpdiblcb = -7.472711488e-7   drout = 0.56   pscbe1 = 7.605327747e+08 wpscbe1 = 4.715364153e+1   pscbe2 = 2.143043264e-08 wpscbe2 = -1.914565709e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -7.056290860e+00 wbeta0 = 1.595161036e-5   agidl = -7.716882287e-10 wagidl = 1.455558301e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = -2.309179502e+00 wegidl = 3.821517620e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.008388520e-01 wkt1 = 7.185448865e-8   kt2 = 6.199812117e-03 wkt2 = -7.004929333e-8   at = 0.0   ute = -9.352406739e-01 wute = 9.605438566e-7   ua1 = 4.573721170e-09 wua1 = -3.290830488e-15   ub1 = -4.640434766e-18 wub1 = 4.694667375e-24   uc1 = 1.759038456e-09 wuc1 = -2.114698604e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.067637354e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.494805350e-07 wvth0 = -5.808470110e-08 pvth0 = -5.256613855e-13   k1 = 4.397755293e-01 lk1 = 1.318007683e-06 wk1 = 1.907573141e-08 pk1 = -1.655626333e-12   k2 = 4.434582590e-02 lk2 = -3.218464608e-07 wk2 = -3.329561876e-08 pk2 = 4.087916660e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.270568712e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.281413302e-07 wvoff = -8.069278040e-08 pvoff = -5.962699552e-13   nfactor = {4.380983004e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.650228724e-06 wnfactor = -2.644512126e-06 pnfactor = -5.862773765e-12   eta0 = 0.08   etab = -0.07   u0 = 1.322690091e-02 lu0 = -7.904715701e-08 wu0 = -3.722084636e-09 pu0 = 9.497179904e-14   ua = 3.818802820e-09 lua = -2.240935839e-14 wua = -5.446732186e-15 pua = 2.705951788e-20   ub = -4.769561350e-18 lub = 1.472146608e-23 wub = 7.347485777e-24 pub = -1.813312030e-29   uc = -3.636248073e-10 luc = 1.123700191e-15 wuc = 3.502476939e-16 puc = -1.353299299e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.014219252e+04 lvsat = 6.452543079e-01 wvsat = 2.252699363e-01 pvsat = -1.813019650e-6   a0 = 2.829046595e+00 la0 = 1.198941678e-06 wa0 = -1.815360532e-06 pa0 = -2.377678204e-12   ags = 9.633594688e-01 lags = -5.554956170e-07 wags = -8.413478230e-07 pags = 8.741891683e-13   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -1.500864350e-01 lketa = 2.315984488e-07 wketa = 1.785450541e-07 pketa = -2.870573172e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -2.852547831e+00 lpclm = 2.144587142e-05 wpclm = 3.700977272e-06 ppclm = -2.662036206e-11   pdiblc1 = 0.39   pdiblc2 = 5.782326522e-03 lpdiblc2 = -4.502275815e-08 wpdiblc2 = -8.601323346e-09 ppdiblc2 = 7.048657094e-14   pdiblcb = 7.649739630e-01 lpdiblcb = -2.377361158e-06 wpdiblcb = -1.214108147e-06 ppdiblcb = 3.756999122e-12   drout = 0.56   pscbe1 = -5.979795625e+08 lpscbe1 = 1.093300162e+04 wpscbe1 = 2.186434312e+03 ppscbe1 = -1.721644950e-2   pscbe2 = 9.013125867e-08 lpscbe2 = -5.528887902e-13 wpscbe2 = -1.284551541e-13 ppscbe2 = 8.796982375e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -1.346157279e+01 lbeta0 = 5.154826779e-05 wbeta0 = 2.018518815e-05 pbeta0 = -3.407088148e-11   agidl = -1.344340505e-09 lagidl = 4.608576675e-15 wagidl = 2.437646410e-15 pagidl = -7.903624130e-21   bgidl = 1.838528210e+08 lbgidl = 6.568168863e+03 wbgidl = 9.763013722e+02 pbgidl = -7.857053776e-3   cgidl = 300.0   egidl = -4.747133641e+00 legidl = 1.962010638e-05 wegidl = 7.688678490e-06 pegidl = -3.112204058e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -8.331366915e-01 lkt1 = 2.674258245e-06 wkt1 = 5.110724838e-07 pkt1 = -3.534727601e-12   kt2 = 2.108599956e-02 lkt2 = -1.198006872e-07 wkt2 = -8.308412010e-08 pkt2 = 1.049013530e-13   at = -4.569739486e+05 lat = 3.677623519e+00 wat = 4.368817946e-01 pat = -3.515926385e-6   ute = 1.193154753e+00 lute = -1.712884750e-05 wute = -1.624569629e-06 pute = 2.080441168e-11   ua1 = 2.011449187e-08 lua1 = -1.250686259e-13 wua1 = -2.338838611e-14 pua1 = 1.617406057e-19   ub1 = -1.989063906e-17 lub1 = 1.227302128e-22 wub1 = 2.479052646e-23 pub1 = -1.617269523e-28   uc1 = 3.271217154e-09 luc1 = -1.216967392e-14 wuc1 = -3.927089793e-15 puc1 = 1.458571651e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-8.347873334e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.930439570e-07 wvth0 = -3.304618941e-07 pvth0 = 5.768602070e-13   k1 = 1.082318791e+00 lk1 = -1.282862868e-06 wk1 = -7.649554533e-07 pk1 = 1.517955496e-12   k2 = -1.034394825e-01 lk2 = 2.763552160e-07 wk2 = 1.485389943e-07 pk2 = -3.272339348e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -3.780797065e-01 ldsub = 3.797135584e-06 wdsub = 1.488012049e-06 pdsub = -6.023137972e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {1.531464368e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.060586149e-07 wvoff = -4.507545624e-07 pvoff = 9.016568743e-13   nfactor = {1.042601980e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.281872011e-05 wnfactor = -1.161185260e-05 pnfactor = 3.043500281e-11   eta0 = -1.696721945e-01 leta0 = 1.010616867e-06 weta0 = 3.960380244e-07 peta0 = -1.603072814e-12   etab = 1.482708089e-01 letab = -8.835111237e-07 wetab = -3.462281418e-07 petab = 1.401453617e-12   u0 = -1.865119852e-02 lu0 = 4.998821693e-08 wu0 = 3.402719341e-08 pu0 = -5.782878492e-14   ua = -3.317735068e-09 lua = 6.477741261e-15 wua = 3.007615175e-15 pua = -7.161778008e-21   ub = -1.414691717e-18 lub = 1.141708656e-24 wub = 3.268875712e-24 pub = -1.623824441e-30   uc = -3.921074885e-11 luc = -1.894549245e-16 wuc = -4.357604685e-17 puc = 2.408105937e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 4.301114354e+05 lvsat = -7.713424441e-01 wvsat = -4.505888169e-01 pvsat = 9.227045146e-7   a0 = 4.978920215e+00 la0 = -7.503263013e-06 wa0 = -4.617269925e-06 pa0 = 8.963820590e-12   ags = 1.618499918e+00 lags = -3.207356749e-06 wags = -1.736439019e-06 pags = 4.497316934e-12   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -1.899744278e-01 lketa = 3.930560688e-07 wketa = 2.352585938e-07 pketa = -5.166209652e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.560810097e+00 lpclm = -1.260950846e-05 wpclm = -7.325662066e-06 ppclm = 1.801299299e-11   pdiblc1 = 0.39   pdiblc2 = -1.035352241e-02 lpdiblc2 = 2.029152775e-08 wpdiblc2 = 1.676412844e-08 ppdiblc2 = -3.218707065e-14   pdiblcb = 3.851378498e-01 lpdiblcb = -8.398700353e-07 wpdiblcb = -5.787187409e-07 ppdiblcb = 1.185085770e-12   drout = 0.56   pscbe1 = 3.412778408e+09 lpscbe1 = -5.301644219e+03 wpscbe1 = -4.144472720e+03 ppscbe1 = 8.409637713e-3   pscbe2 = -7.456430807e-08 lpscbe2 = 1.137618075e-13 wpscbe2 = 1.451323265e-13 ppscbe2 = -2.277223268e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -1.277687840e+01 lbeta0 = 4.877677896e-05 wbeta0 = 2.904306461e-05 pbeta0 = -6.992557238e-11   agidl = -4.237386933e-10 lagidl = 8.821876756e-16 wagidl = 8.307710749e-16 pagidl = -1.399354321e-21   bgidl = 1.575015195e+09 lbgidl = 9.370565834e+02 wbgidl = -6.878515772e+02 pbgidl = -1.120937071e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 8.733558725e-02 lkt1 = -1.051606433e-06 wkt1 = -6.806874897e-07 pkt1 = 1.289248626e-12   kt2 = 2.219120556e-02 lkt2 = -1.242743124e-07 wkt2 = -9.871940278e-08 pkt2 = 1.681894594e-13   at = 8.141329198e+05 lat = -1.467531085e+00 wat = -8.513566346e-01 pat = 1.698572923e-6   ute = -6.362047684e+00 lute = 1.345291204e-05 wute = 7.451230745e-06 pute = -1.593238618e-11   ua1 = -2.387616587e-08 lua1 = 5.299565872e-14 wua1 = 3.254098787e-14 pua1 = -6.464891605e-20   ub1 = 2.191096329e-17 lub1 = -4.647326810e-23 wub1 = -2.961921375e-23 pub1 = 5.851143382e-29   uc1 = 3.219910101e-10 luc1 = -2.318700692e-16 wuc1 = -3.630772034e-16 puc1 = 1.593954456e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.102033643e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.421635515e-08 wvth0 = -2.704415684e-08 pvth0 = -4.447104998e-14   k1 = 6.762255142e-01 lk1 = -4.512752081e-07 wk1 = -3.877424770e-07 pk1 = 7.455081931e-13   k2 = -5.734745954e-02 lk2 = 1.819691237e-07 wk2 = 1.355949202e-07 pk2 = -3.007273835e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.407399387e+00 ldsub = -1.906898868e-06 wdsub = -3.213326664e-06 pdsub = 3.604145911e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.432985506e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.057715191e-07 wvoff = 5.163129301e-08 pvoff = -1.271163207e-13   nfactor = {-3.398211777e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.490195716e-06 wnfactor = 6.893151128e-06 pnfactor = -7.459081193e-12   eta0 = 4.369365558e-01 leta0 = -2.315813666e-07 weta0 = -7.971967195e-07 peta0 = 8.404034634e-13   etab = 3.148499546e-01 letab = -1.224627734e-06 wetab = 6.572928126e-07 petab = -6.535315057e-13   u0 = 7.482636904e-03 lu0 = -3.527997904e-09 wu0 = 4.742323879e-09 pu0 = 2.140038790e-15   ua = -4.214741941e-10 lua = 5.468506501e-16 wua = 4.559605116e-16 pua = -1.936563380e-21   ub = 1.825727964e-19 lub = -2.129129683e-24 wub = 4.301760363e-25 pub = 4.189193787e-30   uc = -2.720506096e-10 luc = 2.873487214e-16 wuc = 2.354599153e-16 puc = -3.305922737e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -2.229677432e+04 lvsat = 1.550877775e-01 wvsat = 9.818934862e-02 pvsat = -2.010696934e-7   a0 = 1.678496825e-01 la0 = 2.348726946e-06 wa0 = 1.507775543e-06 pa0 = -3.578894393e-12   ags = -7.938414224e-02 lags = 2.695277826e-07 wags = 2.782836317e-07 pags = 3.716182579e-13   a1 = 0.0   a2 = 1.442727854e+00 la2 = -1.316162031e-06 wa2 = -1.019515489e-06 pa2 = 2.087738330e-12   b0 = 0.0   b1 = 0.0   keta = 2.380971008e-02 lketa = -4.472574410e-08 wketa = -4.135893673e-08 pketa = 4.982949833e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.285746620e+00 lpclm = 1.410699218e-06 wpclm = 2.077329257e-06 ppclm = -1.242217564e-12   pdiblc1 = -6.570046958e-01 lpdiblc1 = 2.144030041e-06 wpdiblc1 = 1.692397598e-06 ppdiblc1 = -3.465649491e-12   pdiblc2 = -1.360699847e-03 lpdiblc2 = 1.876250532e-09 wpdiblc2 = 2.142092459e-09 ppdiblc2 = -2.244430926e-15   pdiblcb = -0.025   drout = 1.399611601e-01 ldrout = 8.601450355e-07 wdrout = -4.902417129e-08 pdrout = 1.003904724e-13   pscbe1 = 8.047162889e+08 lpscbe1 = 3.908018667e+01 wpscbe1 = -7.481128334e+00 ppscbe1 = -6.199024266e-5   pscbe2 = -4.901717115e-08 lpscbe2 = 6.144701917e-14 wpscbe2 = 7.004169433e-14 ppscbe2 = -7.395360756e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.469911039e+00 lbeta0 = 3.220359710e-06 wbeta0 = -4.341417970e-06 pbeta0 = -1.561663555e-12   agidl = 1.221102050e-09 lagidl = -2.486076077e-15 wagidl = -1.778327947e-15 pagidl = 3.943493428e-21   bgidl = 2.098137327e+09 lbgidl = -1.341798386e+02 wbgidl = -1.313627010e+03 pbgidl = 1.605102167e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.986590275e-01 lkt1 = -5.639881112e-08 wkt1 = -7.133318936e-08 pkt1 = 4.142812361e-14   kt2 = -7.563189251e-02 lkt2 = 7.604538229e-08 wkt2 = 2.306980524e-08 pkt2 = -8.120743606e-14   at = -3.937344349e+04 lat = 2.802579079e-01 wat = 1.636785477e-01 pat = -3.799907473e-7   ute = -2.943706079e+00 lute = 6.452917558e-06 wute = 4.669400781e-06 pute = -1.023582432e-11   ua1 = -7.525841530e-09 lua1 = 1.951387329e-14 wua1 = 1.643753148e-14 pua1 = -3.167266064e-20   ub1 = 7.058656686e-18 lub1 = -1.605908595e-23 wub1 = -1.362688442e-23 pub1 = 2.576274162e-29   uc1 = 1.053225321e-09 luc1 = -1.729273411e-15 wuc1 = -1.416498318e-15 puc1 = 2.316564869e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.081832354e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.304994912e-08 wvth0 = -7.084136737e-08 pvth0 = 1.418572275e-15   k1 = -2.872309938e-01 lk1 = 5.582104345e-07 wk1 = 9.612765546e-07 pk1 = -6.679602228e-13   k2 = 3.471420021e-01 lk2 = -2.418448221e-07 wk2 = -4.469200290e-07 pk2 = 3.096172174e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.342608392e+00 ldsub = 3.070040534e-06 wdsub = 4.405425147e-06 pdsub = -4.378591767e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.433105301e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.006570898e-09 wvoff = -7.061471531e-08 pvoff = 9.699906798e-16   nfactor = {-1.681961476e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.691951557e-06 wnfactor = 5.500111382e-06 pnfactor = -5.999488974e-12   eta0 = 1.757848766e+00 leta0 = -1.615600158e-06 weta0 = -2.193467536e-06 peta0 = 2.303381119e-12   etab = -1.789344850e+00 letab = 9.800949781e-07 wetab = 7.099434879e-08 petab = -3.922263277e-14   u0 = -5.479977332e-03 lu0 = 1.005390523e-08 wu0 = 2.579116343e-08 pu0 = -1.991440907e-14   ua = -1.361428283e-09 lua = 1.531711046e-15 wua = 1.680808748e-15 pua = -3.219928741e-21   ub = -2.419937349e-18 lub = 5.977153843e-25 wub = 5.018039234e-24 pub = -6.178545746e-31   uc = 4.713071834e-11 luc = -4.708149452e-17 wuc = -1.796800838e-16 puc = 1.043810389e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.916768343e+05 lvsat = -4.882184203e-01 wvsat = -8.448281262e-01 pvsat = 7.870004413e-7   a0 = 2.196663909e+00 la0 = 2.229861203e-07 wa0 = -1.524868256e-06 pa0 = -4.013660364e-13   ags = -1.009657450e+00 lags = 1.244244898e-06 wags = 1.341851581e-06 pags = -7.427616506e-13   a1 = 0.0   a2 = -7.378228411e-01 la2 = 9.685644736e-07 wa2 = 2.091801885e-06 pa2 = -1.172222232e-12   b0 = 0.0   b1 = 0.0   keta = 4.295513683e-02 lketa = -6.478584361e-08 wketa = -3.628379702e-08 pketa = 4.451189382e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -2.941610810e+00 lpclm = 3.145672320e-06 wpclm = 5.503052005e-06 ppclm = -4.831604217e-12   pdiblc1 = -1.507649800e+00 lpdiblc1 = 3.035314715e-06 wpdiblc1 = 1.886846503e-06 ppdiblc1 = -3.669388192e-12   pdiblc2 = -3.498168347e-03 lpdiblc2 = 4.115836590e-09 wpdiblc2 = 5.209930638e-09 ppdiblc2 = -5.458835074e-15   pdiblcb = -1.165260703e-01 lpdiblcb = 9.589872833e-08 wpdiblcb = 1.023166877e-07 ppdiblcb = -1.072048675e-13   drout = 1.046251774e+00 ldrout = -8.944361226e-08 wdrout = -5.532785177e-08 pdrout = 1.069953112e-13   pscbe1 = 9.270133664e+08 lpscbe1 = -8.905963369e+01 wpscbe1 = -1.862744543e+02 ppscbe1 = 1.253449345e-4   pscbe2 = 1.036039464e-08 lpscbe2 = -7.673098240e-16 wpscbe2 = -1.614314094e-15 ppscbe2 = 1.125766670e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.433474524e+01 lbeta0 = -1.876891949e-06 wbeta0 = -9.394457301e-06 pbeta0 = 3.732784729e-12   agidl = -2.211760633e-09 lagidl = 1.110791621e-15 wagidl = 3.666988693e-15 pagidl = -1.761973214e-21   bgidl = 2.161044317e+09 lbgidl = -2.000922105e+02 wbgidl = -1.388878365e+03 pbgidl = 2.393567052e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.665921516e-01 lkt1 = 1.195573180e-07 wkt1 = 1.820313701e-07 pkt1 = -2.240409277e-13   kt2 = 9.593964179e-02 lkt2 = -1.037229821e-07 wkt2 = -1.936839481e-07 pkt2 = 1.459017278e-13   at = 4.399683371e+05 lat = -2.219844262e-01 wat = -4.174699692e-01 pat = 2.289221399e-7   ute = 6.159074426e+00 lute = -3.084748285e-06 wute = -9.734965015e-06 pute = 4.856710048e-12   ua1 = 2.229532515e-08 lua1 = -1.173199962e-14 wua1 = -3.111278290e-14 pua1 = 1.814937000e-20   ub1 = -1.806355025e-17 lub1 = 1.026333443e-23 wub1 = 2.704732695e-23 pub1 = -1.685468019e-29   uc1 = -1.594889442e-09 luc1 = 1.045355036e-15 wuc1 = 2.331593588e-15 puc1 = -1.610592128e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.058404233e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.021661023e-08 wvth0 = -1.907579282e-08 pvth0 = -2.693731532e-14   k1 = -1.094633757e+00 lk1 = 1.000485483e-06 wk1 = 1.897777277e-06 pk1 = -1.180951906e-12   k2 = 5.712387404e-01 lk2 = -3.645994129e-07 wk2 = -6.574347281e-07 pk2 = 4.249319067e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 7.397286466e+00 ldsub = -2.265230372e-06 wdsub = -9.320613658e-06 pdsub = 3.140189139e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {5.966693964e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.101794126e-07 wvoff = -3.077063264e-07 pvoff = 1.308428480e-13   nfactor = {8.757451365e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.026497812e-06 wnfactor = -1.244814045e-05 pnfactor = 3.832114673e-12   eta0 = -3.194417199e+00 leta0 = 1.097127332e-06 weta0 = 4.407417755e-06 peta0 = -1.312418822e-12   etab = 2.751398957e-03 letab = -1.570544866e-09 wetab = -4.920571238e-09 petab = 2.361662551e-15   u0 = 2.703692680e-02 lu0 = -7.758041931e-09 wu0 = -2.972772035e-08 pu0 = 1.049744749e-14   ua = 9.661563786e-09 lua = -4.506408435e-15 wua = -1.593538186e-14 pua = 6.429780072e-21   ub = -9.899499218e-18 lub = 4.694832387e-24 wub = 1.620250198e-23 pub = -6.744423655e-30   uc = -4.455541808e-11 luc = 3.141878852e-18 wuc = -2.469106035e-17 puc = 1.948192653e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -9.136143481e+05 lvsat = 3.363424571e-01 wvsat = 1.523275358e+00 pvsat = -5.101874447e-7   a0 = 4.199268355e+00 la0 = -8.739905299e-07 wa0 = -3.990400904e-06 pa0 = 9.491911100e-13   ags = 2.290032349e+00 lags = -5.632426820e-07 wags = -1.639653323e-06 pags = 8.904321982e-13   a1 = 0.0   a2 = 1.969040982e+00 la2 = -5.141878572e-07 wa2 = -9.002067655e-07 pa2 = 4.667253071e-13   b0 = 0.0   b1 = 0.0   keta = 6.717458365e-02 lketa = -7.805265109e-08 wketa = -1.317536746e-07 pketa = 9.680790603e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.911112549e+00 lpclm = -1.155853218e-06 wpclm = -6.711716245e-06 ppclm = 1.859340461e-12   pdiblc1 = 8.095425594e+00 lpdiblc1 = -2.225009909e-06 wpdiblc1 = -1.023763918e-05 ppdiblc1 = 2.972101951e-12   pdiblc2 = -5.475130596e-03 lpdiblc2 = 5.198767086e-09 wpdiblc2 = -6.444337316e-09 ppdiblc2 = 9.250815544e-16   pdiblcb = 4.255137896e-01 lpdiblcb = -2.010171559e-07 wpdiblcb = -2.517423099e-07 ppdiblcb = 8.673979996e-14   drout = 4.057755920e-01 ldrout = 2.613932282e-07 wdrout = 1.438826016e-06 pdrout = -7.114648237e-13   pscbe1 = 7.219546834e+08 lpscbe1 = 2.326638638e+01 wpscbe1 = 9.340155409e+01 ppscbe1 = -2.785459102e-5   pscbe2 = 7.927231228e-09 lpscbe2 = 5.655162622e-16 wpscbe2 = 1.922694804e-15 ppscbe2 = -8.117183789e-22   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.328281730e+01 lbeta0 = -1.300672117e-06 wbeta0 = -5.712659906e-06 pbeta0 = 1.715988161e-12   agidl = -1.590590223e-09 lagidl = 7.705299991e-16 wagidl = 2.264969698e-15 pagidl = -9.939822589e-22   bgidl = 3.694827528e+09 lbgidl = -1.040260309e+03 wbgidl = -3.594619423e+03 pbgidl = 1.447606513e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.543401000e-01 lkt1 = -1.062640495e-07 wkt1 = -4.884731688e-07 pkt1 = 1.432446961e-13   kt2 = -1.618759906e-01 lkt2 = 3.750197598e-08 wkt2 = 1.835168749e-07 pkt2 = -6.071945297e-14   at = 2.915150971e+05 lat = -1.406654527e-01 wat = -3.594135636e-01 pat = 1.971202924e-7   ute = -1.903942124e+00 lute = 1.331970605e-06 wute = 2.988369281e-06 pute = -2.112814397e-12   ua1 = -1.149906650e-09 lua1 = 1.110712225e-15 wua1 = 7.688718866e-15 pua1 = -3.105122624e-21   ub1 = 3.111467768e-18 lub1 = -1.335811067e-24 wub1 = -9.865868300e-24 pub1 = 3.365445336e-30   uc1 = 4.354003413e-10 luc1 = -6.678695053e-17 wuc1 = -8.851272981e-16 puc1 = 1.514471555e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-8.070513571e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.774882328e-08 wvth0 = -4.005489098e-07 pvth0 = 9.160303144e-14   k1 = 8.088631369e+00 lk1 = -1.833058996e-06 wk1 = -1.130539765e-05 pk1 = 2.907656837e-12   k2 = -2.800423071e+00 lk2 = 6.759004225e-07 wk2 = 4.175624391e-06 pk2 = -1.072134879e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.099452272e+00 ldsub = 1.539108370e-06 wdsub = 8.980858031e-06 pdsub = -2.441382948e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-7.680717429e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.440818792e-07 wvoff = 8.577609587e-07 pvoff = -2.285472874e-13   nfactor = {-8.756330217e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.370709853e-06 wnfactor = 1.740689333e-05 pnfactor = -5.346727832e-12   eta0 = -3.016567052e+00 leta0 = 1.103779644e-06 weta0 = 5.562228868e-06 peta0 = -1.750850592e-12   etab = -2.884269014e-01 letab = 8.999544209e-08 wetab = 4.565205856e-07 petab = -1.427536501e-13   u0 = -2.375343623e-02 lu0 = 7.786587317e-09 wu0 = 4.476384230e-08 pu0 = -1.235133397e-14   ua = -2.007570721e-08 lua = 4.596869804e-15 wua = 2.882217113e-14 pua = -7.291701983e-21   ub = 2.094491888e-17 lub = -4.746190942e-24 wub = -3.036416730e-23 pub = 7.528559950e-30   uc = -2.106014483e-10 luc = 5.558838815e-17 wuc = 3.208580826e-16 puc = -8.817608011e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 4.377872415e+05 lvsat = -6.984315883e-02 wvsat = -5.420142702e-01 pvsat = 1.107874535e-7   a0 = 1.969725246e+00 la0 = -2.220822914e-07 wa0 = -1.921918739e-06 pa0 = 3.522740373e-13   ags = -2.578886351e+00 lags = 9.372156294e-07 wags = 6.073502011e-06 pags = -1.486641422e-12   a1 = 0.0   a2 = -1.355374553e+00 la2 = 5.029000147e-07 wa2 = 3.201411186e-06 pa2 = -7.977160961e-13   b0 = 0.0   b1 = 0.0   keta = -3.474194822e-01 lketa = 4.799516350e-08 wketa = 4.352104800e-07 pketa = -7.613146419e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.924519023e+00 lpclm = -2.817359987e-07 wpclm = -1.887344204e-06 ppclm = 4.468986567e-13   pdiblc1 = 3.618275295e-01 lpdiblc1 = 8.230741771e-08 wpdiblc1 = 1.581615172e-07 ppdiblc1 = -1.305586598e-13   pdiblc2 = -2.345200644e-03 lpdiblc2 = 4.510341439e-09 wpdiblc2 = 1.939107674e-08 ppdiblc2 = -7.154447921e-15   pdiblcb = -3.408533497e-01 lpdiblcb = 2.873997386e-08 wpdiblcb = 1.843788837e-07 ppdiblcb = -4.558826622e-14   drout = 2.809766946e+00 ldrout = -4.804001886e-07 wdrout = -3.371303641e-06 pdrout = 7.620261519e-13   pscbe1 = 8.003993042e+08 lpscbe1 = -9.773916597e-02 wpscbe1 = -6.333882571e-01 ppscbe1 = 1.550369927e-7   pscbe2 = 1.064539244e-08 lpscbe2 = -2.578075603e-16 wpscbe2 = -2.102409006e-15 ppscbe2 = 4.089426019e-22   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.312786762e+00 lbeta0 = 1.763388763e-06 wbeta0 = 8.936209141e-06 pbeta0 = -2.797143684e-12   agidl = 1.759831459e-08 lagidl = -5.225667892e-15 wagidl = -2.740654304e-14 pagidl = 8.289121631e-21   bgidl = -2.591207123e+09 lbgidl = 8.790376992e+02 wbgidl = 5.696487619e+03 pbgidl = -1.394357728e-3   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -8.005149003e-01 lkt1 = 9.106899963e-08 wkt1 = 4.514969984e-07 pkt1 = -1.444565614e-13   kt2 = -3.762382566e-02 lkt2 = 5.314917424e-10 wkt2 = -1.771531472e-08 pkt2 = -8.430692095e-16   at = -6.398344561e+05 lat = 1.444695003e-01 wat = 1.030582627e+00 pat = -2.291621443e-7   ute = 8.844867161e+00 lute = -1.975443522e-06 wute = -1.406173596e-05 pute = 3.133511729e-12   ua1 = 4.083339950e-09 lua1 = -4.731723182e-16 wua1 = -5.123465743e-15 pua1 = 7.505610726e-22   ub1 = -1.028797524e-18 lub1 = -1.088206267e-25 wub1 = 8.877307322e-25 pub1 = 1.726147603e-31   uc1 = 7.609033716e-10 luc1 = -1.730600395e-16 wuc1 = -1.248625308e-15 puc1 = 2.745133726e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-9.530712863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.200679512e-08 wvth0 = -1.338639995e-07 pvth0 = 2.632523254e-14   k1 = -3.109488982e+00 lk1 = 9.079609132e-07 wk1 = 5.010765097e-06 pk1 = -1.086131899e-12   k2 = 1.390786837e+00 lk2 = -3.500029827e-07 wk2 = -1.914947142e-06 pk2 = 4.186847680e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.946356194e+00 ldsub = -1.898954397e-06 wdsub = -1.027344884e-05 pdsub = 2.271590017e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-4.314517267e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.168571476e-08 wvoff = 2.255196698e-07 pvoff = -7.379042594e-14   nfactor = {5.896805875e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.160115334e-07 wnfactor = -5.492208872e-06 pnfactor = 2.583999087e-13   eta0 = 1.132807652e+01 leta0 = -2.407430486e-06 weta0 = -1.335594487e-05 peta0 = 2.879845385e-12   etab = 1.383463998e+00 letab = -3.192416528e-07 wetab = -1.686838544e-06 petab = 3.818870808e-13   u0 = 8.223753074e-03 lu0 = -4.062919389e-11 wu0 = -5.894664141e-09 pu0 = 4.860194186e-17   ua = -5.300583552e-09 lua = 9.802889100e-16 wua = 3.823502886e-15 pua = -1.172652963e-21   ub = 8.028119405e-18 lub = -1.584481349e-24 wub = -7.350572546e-24 pub = 1.895407293e-30   uc = 1.186221205e-10 luc = -2.499731090e-17 wuc = -1.615386627e-16 puc = 2.990258321e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.255244451e+06 lvsat = -2.699362474e-01 wvsat = -1.408601640e+00 pvsat = 3.229063771e-7   a0 = 4.109653868e+00 la0 = -7.458833199e-07 wa0 = -4.127926126e-06 pa0 = 8.922494956e-13   ags = 1.249999095e+00 lags = 1.944347687e-13 wags = 1.082943044e-12 pags = -2.325890929e-19   a1 = 0.0   a2 = -3.431427501e-01 la2 = 2.551309750e-07 wa2 = 1.189276533e-06 pa2 = -3.051958365e-13   b0 = -6.136079655e-23 lb0 = 1.501958897e-29 wb0 = 7.340174837e-29 pb0 = -1.796691296e-35   b1 = 0.0   keta = -1.761694040e+00 lketa = 3.941742184e-07 wketa = 2.050540270e-06 pketa = -4.715238136e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.756449969e+00 lpclm = -4.853718962e-07 wpclm = -2.433636666e-06 ppclm = 5.806173941e-13   pdiblc1 = 9.301381160e+00 lpdiblc1 = -2.105871822e-06 wpdiblc1 = -1.066675901e-05 ppdiblc1 = 2.519111261e-12   pdiblc2 = 1.870125856e-01 lpdiblc2 = -4.183971069e-08 wpdiblc2 = -2.143110935e-07 ppdiblc2 = 5.005000080e-14   pdiblcb = -4.579998106e+00 lpdiblcb = 1.066376632e-06 wpdiblcb = 5.209588095e-06 ppdiblcb = -1.275633851e-12   drout = -8.342162613e+00 ldrout = 2.249313369e-06 wdrout = 1.073441296e-05 pdrout = -2.690700630e-12   pscbe1 = 8.108769046e+08 lpscbe1 = -2.662393817e+00 wpscbe1 = -1.301130139e+01 ppscbe1 = 3.184840681e-6   pscbe2 = 5.487314447e-08 lpscbe2 = -1.108365556e-14 wpscbe2 = -5.459829649e-14 ppscbe2 = 1.325862346e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.064814829e+01 lbeta0 = -4.927624356e-06 wbeta0 = -2.657283231e-05 pbeta0 = 5.894581938e-12   agidl = -1.394089428e-08 lagidl = 2.494341961e-15 wagidl = 1.864772437e-14 pagidl = -2.983811673e-21   bgidl = 9.999991834e+08 lbgidl = 1.753835487e-04 wbgidl = 9.768334961e-04 pbgidl = -2.097994127e-10   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 4.014059267e-01 lkt1 = -2.031311708e-07 wkt1 = -1.131379391e-06 pkt1 = 2.429920067e-13   kt2 = 9.118267863e-02 lkt2 = -3.099712034e-08 wkt2 = -1.726446027e-07 pkt2 = 3.707974726e-14   at = -6.143862522e+05 lat = 1.382404161e-01 wat = 7.699574209e-01 pat = -1.653676095e-7   ute = 8.316034960e+00 lute = -1.845998620e-06 wute = -1.028165586e-05 pute = 2.208242621e-12   ua1 = 1.308151569e-08 lua1 = -2.675700784e-15 wua1 = -1.513346606e-14 pua1 = 3.200758900e-21   ub1 = -1.100667358e-17 lub1 = 2.333513986e-24 wub1 = 1.299696927e-23 pub1 = -2.791424102e-30   uc1 = 8.147454870e-10 luc1 = -1.862392433e-16 wuc1 = -1.037296414e-15 puc1 = 2.227853425e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-6.811440510e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.696743820e-06 wvth0 = -4.809829691e-07 pvth0 = 9.642638342e-12   k1 = 1.007111856e+00 lk1 = -1.121861794e-05 wk1 = -6.120138164e-07 pk1 = 1.226951529e-11   k2 = -2.299981727e-01 lk2 = 4.991520735e-06 wk2 = 2.924584984e-07 pk2 = -5.863142172e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.012882948e-04 lcit = -1.830127195e-09 wcit = -1.092019795e-10 pcit = 2.189256714e-15   voff = {-5.141530527e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.043946193e-06 wvoff = -1.340365889e-07 pvoff = 2.687135375e-12   nfactor = {9.646444605e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.579785060e-04 wnfactor = -8.389300854e-06 pnfactor = 1.681868159e-10   eta0 = 0.08   etab = -0.07   u0 = 1.408832780e-02 lu0 = -7.878831307e-08 wu0 = -7.185321429e-09 pu0 = 1.440497073e-13   ua = 3.975471886e-09 lua = -9.389692028e-14 wua = -4.961841022e-15 pua = 9.947387239e-20   ub = -3.170403471e-18 lub = 8.998894044e-23 wub = 3.803165665e-24 pub = -7.624500953e-29   uc = -1.519758743e-10 luc = 1.607810812e-15 wuc = 3.994788540e-17 puc = -8.008662182e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.166015950e+05 lvsat = -1.516196373e+01 wvsat = -9.046964672e-01 pvsat = 1.813715122e-5   a0 = 3.485692867e+00 la0 = -4.555283235e-05 wa0 = -2.069066605e-06 pa0 = 4.148018175e-11   ags = 3.481073890e+00 lags = -6.413814269e-05 wags = -3.601766201e-06 pags = 7.220739839e-11   a1 = 0.0   a2 = -8.039752190e-01 la2 = 3.215613430e-05 wa2 = 1.918726484e-06 pa2 = -3.846619684e-11   b0 = -2.587306380e-07 lb0 = 5.186973616e-12 wb0 = 3.095018685e-13 pb0 = -6.204823822e-18   b1 = 3.773587581e-08 lb1 = -7.565203477e-13 wb1 = -4.514086220e-14 pb1 = 9.049738486e-19   keta = -5.537279577e-01 lketa = 1.106352016e-05 wketa = 6.162185814e-07 pketa = -1.235381147e-11   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.658554649e-01 lpclm = -6.513451628e-06 wpclm = -5.095478967e-07 ppclm = 1.021530159e-11   pdiblc1 = 0.39   pdiblc2 = -9.063500624e-03 lpdiblc2 = 1.881042361e-07 wpdiblc2 = 1.117567037e-08 ppdiblc2 = -2.240473252e-13   pdiblcb = 2.145428258e+00 lpdiblcb = -4.612086443e-05 wpdiblcb = -2.522218755e-06 ppdiblcb = 5.056487411e-11   drout = 0.56   pscbe1 = 6.959287808e+08 lpscbe1 = 2.085419057e+03 wpscbe1 = 1.099362556e+02 ppscbe1 = -2.203977316e-3   pscbe2 = 3.741205363e-09 lpscbe2 = 3.376561414e-14 wpscbe2 = 7.901648617e-15 ppscbe2 = -1.584104736e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.043514835e-09 lalpha0 = -1.891537311e-14 walpha0 = -1.128662638e-15 palpha0 = 2.262717461e-20   alpha1 = 1.043514835e-09 lalpha1 = -1.891537311e-14 walpha1 = -1.128662638e-15 palpha1 = 2.262717461e-20   beta0 = -2.525706106e+02 lbeta0 = 5.189350519e-03 wbeta0 = 3.047389122e-04 pbeta0 = -6.109337145e-9   agidl = -1.648136030e-08 lagidl = 3.393378222e-13 wagidl = 1.980041725e-14 pagidl = -3.969543100e-19   bgidl = 1000000000.0   cgidl = 300.0   egidl = -9.683147321e-02 legidl = 1.969255094e-05 pegidl = -1.421085472e-26   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -6.223746595e-01 lkt1 = 3.640739281e-06 wkt1 = 1.951457701e-07 pkt1 = -3.912238490e-12   kt2 = 1.598694947e-01 lkt2 = -4.254698525e-06 wkt2 = -2.323352040e-07 pkt2 = 4.657803894e-12   at = -6.698011811e+05 lat = 1.342802337e+01 wat = 8.012376065e-01 pat = -1.606303126e-5   ute = -2.706909318e+00 lute = 5.161586753e-05 wute = 2.784523594e-06 pute = -5.582350248e-11   ua1 = 6.526630007e-09 lua1 = -9.430284324e-14 wua1 = -4.615101526e-15 pua1 = 9.252251699e-20   ub1 = -6.186347551e-18 lub1 = 1.096705246e-22 wub1 = 5.100426460e-24 pub1 = -1.022522021e-28   uc1 = 4.834104492e-09 luc1 = -9.708868319e-14 wuc1 = -5.142965755e-15 puc1 = 1.031050203e-19   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.114945+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.44751769   k2 = 0.01898311   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.20324992+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7663429+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.0101583   ua = -7.0818604e-10   ub = 1.31832111e-18   uc = -7.1776909e-11   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160310.0   a0 = 1.213479   ags = 0.281809   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -0.0018702   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.14095898   pdiblc1 = 0.39   pdiblc2 = 0.00031929802   pdiblcb = -0.15511953   drout = 0.56   pscbe1 = 799951250.0   pscbe2 = 5.4254628e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.2785893   agidl = 4.4509773e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.88544965   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.4407715   kt2 = -0.052358472   at = 0.0   ute = -0.13226612   ua1 = 1.8227243e-9   ub1 = -7.1588888e-19   uc1 = -8.7612717e-12   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539358e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584525e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-08 wpdiblc2 = -8.673617380e-25 ppdiblc2 = 3.469446952e-30   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 wpscbe2 = -1.323488980e-29 ppscbe2 = 5.293955920e-35   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-7   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23 pub1 = -6.162975822e-45   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308607e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = -1.387778781e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = 2.220446049e-22 ppclm = -1.332267630e-27   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343241e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 wuc1 = -1.292469707e-32 puc1 = -2.584939414e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-08 wk2 = -5.551115123e-23   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = -6.591949209e-23 peta0 = -4.354155925e-28   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = -2.151057110e-22 petab = 8.673617380e-30   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493534e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554778e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463398e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = -2.220446049e-22   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15 pua1 = 6.617444900e-36   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 wuc1 = 1.033975766e-31 puc1 = -2.067951531e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.68 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.141052779e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.423581630e-8   k1 = 5.163560651e-01 lk1 = -1.764191989e-10   k2 = -2.646447971e-02 lk2 = 1.698224276e-08 pk2 = -1.387778781e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.340143070e+00 ldsub = -5.902793436e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.023414834e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.817442602e-9   nfactor = {2.915901967e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.323370700e-6   eta0 = -7.579850000e-02 leta0 = 3.099302733e-7   etab = -1.729996539e+00 letab = 9.473064950e-7   u0 = 1.608035831e-02 lu0 = -6.593709171e-9   ua = 4.365764318e-11 lua = -1.160014925e-15   ub = 1.774933909e-18 lub = 8.121476016e-26   uc = -1.030743287e-10 luc = 4.017669524e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.145642010e+05 lvsat = 1.696810852e-1   a0 = 9.219377220e-01 la0 = -1.125391259e-7   ags = 1.120744390e-01 lags = 6.233271742e-7   a1 = 0.0   a2 = 1.010836186e+00 la2 = -1.136436256e-8   b0 = 0.0   b1 = 0.0   keta = 1.262339765e-02 lketa = -2.757575910e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.658710871e+00 lpclm = -8.933470478e-7   pdiblc1 = 6.967508558e-02 lpdiblc1 = -3.214058779e-8   pdiblc2 = 8.571161110e-04 lpdiblc2 = -4.475215832e-10   pdiblcb = -3.099359191e-02 lpdiblcb = 6.279935762e-9   drout = 1.0   pscbe1 = 7.712957009e+08 lpscbe1 = 1.572349742e+1   pscbe2 = 9.010895465e-09 lpscbe2 = 1.737841029e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.481371233e+00 lbeta0 = 1.243560211e-6   agidl = 8.536887886e-10 lagidl = -3.621444101e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.144215274e-01 lkt1 = -6.773154207e-8   kt2 = -6.597205099e-02 lkt2 = 1.824476986e-08 wkt2 = -1.110223025e-22   at = 9.098087549e+04 lat = -3.061507655e-2   ute = -1.978949816e+00 lute = 9.752585094e-7   ua1 = -3.713662156e-09 lua1 = 3.440115825e-15 wua1 = 1.654361225e-30 pua1 = 8.271806126e-37   ub1 = 4.546885644e-18 lub1 = -3.826474399e-24 pub1 = -1.540743956e-45   uc1 = 3.542254351e-10 luc1 = -3.010327285e-16 wuc1 = -2.067951531e-31   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.69 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.074350799e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.301860543e-9   k1 = 4.918287993e-01 lk1 = 1.325900381e-8   k2 = 2.165076081e-02 lk2 = -9.374083109e-09 pk2 = -6.938893904e-30   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -3.943573436e-01 ldsub = 3.598366204e-07 pdsub = 2.220446049e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.975627001e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.002553889e-10   nfactor = {-1.648674244e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.176990034e-06 pnfactor = -4.440892099e-28   eta0 = 0.49   etab = -1.361993125e-03 letab = 4.037064090e-10   u0 = 2.185793948e-03 lu0 = 1.017385823e-9   ua = -3.659750026e-09 lua = 8.686192116e-16   ub = 3.645115856e-18 lub = -9.432241560e-25 pub = 1.540743956e-45   uc = -6.519611348e-11 luc = 1.942795591e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.597802425e+05 lvsat = -9.015294234e-02 wvsat = 4.656612873e-16   a0 = 8.634598290e-01 la0 = -8.050639808e-8   ags = 9.193506400e-01 lags = 1.811214532e-7   a1 = 0.0   a2 = 1.216505717e+00 la2 = -1.240249899e-7   b0 = 0.0   b1 = 0.0   keta = -4.296598660e-02 lketa = 2.874715860e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.996019656e-01 lpclm = 3.984777661e-07 wpclm = -2.220446049e-22 ppclm = 1.942890293e-28   pdiblc1 = -4.628132577e-01 lpdiblc1 = 2.595432144e-07 wpdiblc1 = -4.163336342e-22 ppdiblc1 = 1.942890293e-28   pdiblc2 = -1.086232749e-02 lpdiblc2 = 5.972096636e-09 wpdiblc2 = 5.421010862e-24 ppdiblc2 = -1.870248748e-30   pdiblcb = 2.150677307e-01 lpdiblcb = -1.285063052e-07 ppdiblcb = 6.938893904e-29   drout = 1.608574059e+00 ldrout = -3.333616552e-7   pscbe1 = 8.000344823e+08 lpscbe1 = -1.888856653e-2   pscbe2 = 9.534523798e-09 lpscbe2 = -1.130464069e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.507272163e+00 lbeta0 = 1.338223295e-7   agidl = 3.028298641e-10 lagidl = -6.039766277e-17   bgidl = 6.898757943e+08 lbgidl = 1.698782868e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.626832716e-01 lkt1 = 1.348253482e-8   kt2 = -8.463546509e-03 lkt2 = -1.325695119e-8   at = -8.939633778e+03 lat = 2.411888042e-2   ute = 5.942098076e-01 lute = -4.342540036e-7   ua1 = 5.277541258e-09 lua1 = -1.485040625e-15   ub1 = -5.135986154e-18 lub1 = 1.477560701e-24   uc1 = -3.045291189e-10 luc1 = 5.981654738e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.70 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-8.869436912e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.810701213e-08 wvth0 = -3.000099100e-07 pvth0 = 8.933545095e-14   k1 = -4.549981676e+00 lk1 = 1.514584118e-06 wk1 = 3.971048753e-06 pk1 = -1.182479042e-12   k2 = 2.018059518e+00 lk2 = -6.038547008e-07 wk2 = -1.646559284e-06 pk2 = 4.903041907e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.805364707e+01 ldsub = -5.133517894e-06 wdsub = -1.884805916e-05 pdsub = 5.612480817e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {9.493163223e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.423121563e-07 wvoff = -1.209031715e-06 pvoff = 3.600194188e-13   nfactor = {1.243458159e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.016651471e-06 wnfactor = -8.232399969e-06 pnfactor = 2.451402901e-12   eta0 = 7.559820324e+00 leta0 = -2.105215747e-06 weta0 = -7.184563379e-06 peta0 = 2.139383360e-12   etab = 7.411262350e-01 letab = -2.206907257e-07 wetab = -7.828078469e-07 petab = 2.331006066e-13   u0 = -1.456630516e-02 lu0 = 6.005742134e-09 wu0 = 3.310387345e-08 pu0 = -9.857505916e-15   ua = -4.312115916e-09 lua = 1.062877464e-15 wua = 9.569702365e-15 pua = -2.849618122e-21   ub = -8.988256999e-19 lub = 4.098480407e-25 wub = -3.825575663e-24 pub = 1.139160793e-30   uc = 2.153333247e-10 luc = -6.410669755e-17 wuc = -1.934420525e-16 puc = 5.760220719e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.538911433e+06 lvsat = -4.412687326e-01 wvsat = -1.853204324e+00 pvsat = 5.518379177e-7   a0 = 6.681110101e+00 la0 = -1.812857208e-06 wa0 = -7.538718089e-06 pa0 = 2.244841779e-12   ags = 2.430890571e+00 lags = -2.689773499e-7   a1 = 0.0   a2 = -7.164474946e-01 la2 = 4.515601527e-07 wa2 = 2.393832108e-06 pa2 = -7.128233560e-13   b0 = 0.0   b1 = 0.0   keta = -6.980987743e-02 lketa = 1.086815545e-08 wketa = 9.899504763e-08 pketa = -2.947825031e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.756023188e-01 lpclm = 3.615537713e-07 wpclm = 1.127624073e-06 ppclm = -3.357782582e-13   pdiblc1 = 8.288488259e-01 lpdiblc1 = -1.250814625e-07 wpdiblc1 = -4.075867799e-07 ppdiblc1 = 1.213691534e-13   pdiblc2 = 6.462168683e-02 lpdiblc2 = -1.650515573e-08 wpdiblc2 = -6.110496773e-08 ppdiblc2 = 1.819553177e-14   pdiblcb = 2.053897663e+00 lpdiblcb = -6.760638882e-07 wpdiblcb = -2.682771958e-06 ppdiblcb = 7.988624197e-13   drout = -3.454820018e+00 ldrout = 1.174390516e-06 wdrout = 4.163933746e-06 pdrout = -1.239915371e-12   pscbe1 = 7.998768488e+08 lpscbe1 = 2.805077190e-2   pscbe2 = -5.429373160e-08 lpscbe2 = 1.889341235e-14 wpscbe2 = 7.560203333e-14 ppscbe2 = -2.251239547e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.083377528e+01 lbeta0 = -6.514452136e-06 wbeta0 = -2.413701598e-05 pbeta0 = 7.187399932e-12   agidl = -3.987398407e-08 lagidl = 1.190325311e-14 wagidl = 4.179332365e-14 pagidl = -1.244500695e-20   bgidl = 2.107586449e+09 lbgidl = -2.522805034e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -2.823373059e-01 lkt1 = -6.999748510e-08 wkt1 = -1.762000254e-07 pkt1 = 5.246796258e-14   kt2 = 1.963604911e-01 lkt2 = -7.424842899e-08 wkt2 = -2.976605763e-07 pkt2 = 8.863587811e-14   at = 7.494182856e+05 lat = -2.017011490e-01 wat = -6.437174263e-01 pat = 1.916829566e-7   ute = -1.999663052e+00 lute = 3.381364872e-07 wute = -9.191767994e-07 pute = 2.737078714e-13   ua1 = -5.958281882e-09 lua1 = 1.860706610e-15 wua1 = 6.929359667e-15 pua1 = -2.063390075e-21   ub1 = 1.224447595e-17 lub1 = -3.697906403e-24 wub1 = -1.498081983e-23 pub1 = 4.460913625e-30   uc1 = 1.527345733e-10 luc1 = -7.634514857e-17 wuc1 = -5.062226731e-16 puc1 = 1.507404565e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.71 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.12e-06 wmax = 1.26e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-2.014599089e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.135780178e-07 wvth0 = 1.135969527e-06 pvth0 = -2.554888594e-13   k1 = 9.333858681e+00 lk1 = -1.770791834e-06 wk1 = -9.874365565e-06 pk1 = 2.118277857e-12   k2 = -3.875890914e+00 lk2 = 7.937682865e-07 wk2 = 4.385221317e-06 pk2 = -9.495310249e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -4.215450277e+01 ldsub = 9.220791585e-06 wdsub = 5.085503388e-05 pdsub = -1.103020596e-11   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.870615409e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.671631460e-07 wvoff = 3.143325319e-06 pvoff = -6.784587045e-13   nfactor = {9.217409714e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.237438625e-07 wnfactor = 4.591229672e-07 pnfactor = 5.068959681e-13   eta0 = -1.279975273e+01 leta0 = 2.721175851e-06 weta0 = 1.550653657e-05 peta0 = -3.255157631e-12   etab = -8.523791594e-01 letab = 1.528882924e-07 wetab = 9.877485880e-07 petab = -1.828898678e-13   u0 = 7.641740268e-02 lu0 = -1.581655605e-08 wu0 = -8.747009000e-08 pu0 = 1.892027047e-14   ua = 2.214238454e-08 lua = -5.333194965e-15 wua = -2.900465372e-14 pua = 6.379738480e-21   ub = -1.448173269e-17 lub = 3.765193130e-24 wub = 1.957643284e-23 pub = -4.504044509e-30   uc = 4.657270967e-10 luc = -1.301814401e-16 wuc = -5.767567426e-16 puc = 1.557272044e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -3.891017945e+06 lvsat = 8.549081140e-01 wvsat = 4.747522118e+00 pvsat = -1.022668443e-6   a0 = -1.211965555e+00 la0 = -1.613231427e-08 wa0 = 2.237965320e-06 pa0 = 1.929799057e-14   ags = 1.25   a1 = 0.0   a2 = 1.406595875e+01 la2 = -3.133101119e-06 wa2 = -1.604735178e-05 pa2 = 3.747915818e-12   b0 = 0.0   b1 = 0.0   keta = 2.698871235e+00 lketa = -6.660246185e-07 wketa = -3.285330650e-06 pketa = 7.967199614e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -2.304966284e+00 lpclm = 8.118434221e-07 wpclm = 3.620991422e-06 ppclm = -9.711530805e-13   pdiblc1 = -1.296299609e+01 lpdiblc1 = 3.241481915e-06 wpdiblc1 = 1.596660152e-05 ppdiblc1 = -3.877564394e-12   pdiblc2 = -3.915340420e-01 lpdiblc2 = 9.391849956e-08 wpdiblc2 = 4.777648959e-07 ppdiblc2 = -1.123483146e-13   pdiblcb = -1.192484680e+01 lpdiblcb = 2.695125220e-06 wpdiblcb = 1.399573113e-05 ppdiblcb = -3.223995032e-12   drout = 2.927086319e+01 ldrout = -6.748387889e-06 wdrout = -3.425949212e-05 pdrout = 8.072637541e-12   pscbe1 = 800000000.0   pscbe2 = 1.194412916e-07 lpscbe2 = -2.222246705e-14 wpscbe2 = -1.318367802e-13 ppscbe2 = 2.658322620e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -5.322814280e+01 lbeta0 = 1.357559736e-05 wbeta0 = 7.376267113e-05 pbeta0 = -1.623956398e-11   agidl = 2.922097509e-08 lagidl = -4.121065554e-15 wagidl = -3.298388496e-14 pagidl = 4.929750490e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -2.096052862e+00 lkt1 = 3.687304740e-07 wkt1 = 1.856160731e-06 pkt1 = -4.410871923e-13   kt2 = -3.005988644e+00 lkt2 = 7.040650448e-07 wkt2 = 3.532290843e-06 pkt2 = -8.422251367e-13   at = -1.698528117e+06 lat = 3.824409550e-01 wat = 2.066842612e+00 pat = -4.574881085e-7   ute = 1.259367067e+01 lute = -3.208709939e-06 wute = -1.539870058e-05 pute = 3.838361508e-12   ua1 = 3.186194956e-08 lua1 = -7.257866598e-15 wua1 = -3.759922203e-14 pua1 = 8.682092276e-21   ub1 = -4.941377573e-17 lub1 = 1.111849870e-23 wub1 = 5.894077389e-23 pub1 = -1.330030394e-29   uc1 = 5.312794375e-10 luc1 = -1.747014922e-16 wuc1 = -6.982052547e-16 puc1 = 2.089835154e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.72 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.136520303e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.325368137e-07 wvth0 = -1.776356839e-21   k1 = 4.276806174e-01 lk1 = 3.976891689e-7   k2 = 4.689033131e-02 lk2 = -5.594776937e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -2.099956519e-06 lcit = 2.425772058e-10 pcit = -9.486769009e-32   voff = {-1.783160135e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.998693471e-7   nfactor = {1.703775898e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.254329181e-6   eta0 = 0.08   etab = -0.07   u0 = 7.285540695e-03 lu0 = 5.759243218e-8   ua = -7.222091363e-10 lua = 2.811318801e-16   ub = 4.302881048e-19 lub = 1.780308588e-23   uc = -1.141547466e-10 luc = 8.495813531e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.006963303e+04 lvsat = 2.009596323e+0   a0 = 1.526779858e+00 la0 = -6.280985109e-06 wa0 = -1.776356839e-21   ags = 7.105961256e-02 lags = 4.225056301e-06 pags = 3.552713679e-27   a1 = 0.0   a2 = 1.012601522e+00 la2 = -4.262187475e-6   b0 = 3.429387608e-08 lb0 = -6.875159114e-13   b1 = -5.001763451e-09 lb1 = 1.002742283e-13   keta = 2.968419166e-02 lketa = -6.325953443e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.656496613e-02 lpclm = 3.158004629e-06 ppclm = 1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 1.517196017e-03 lpdiblc2 = -2.401518953e-8   pdiblcb = -2.425118492e-01 lpdiblcb = 1.752021553e-6   drout = 0.56   pscbe1 = 8.000122166e+08 lpscbe1 = -1.222244938e+0   pscbe2 = 1.122218361e-08 lpscbe2 = -1.162113546e-13   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -2.505971875e-11 lalpha0 = 2.507169103e-15   alpha1 = -2.505971875e-11 lalpha1 = 2.507169103e-15   beta0 = 3.594451880e+01 lbeta0 = -5.947358799e-4   agidl = 2.264916321e-09 lagidl = -3.648331365e-14 pagidl = 5.293955920e-35   bgidl = 1000000000.0   cgidl = 300.0   egidl = -9.683147321e-02 legidl = 1.969255094e-5   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.376181192e-01 lkt1 = -6.321826893e-8   kt2 = -6.009657711e-02 lkt2 = 1.551317903e-7   at = 8.877989434e+04 lat = -1.779839346e+0   ute = -7.062903695e-02 lute = -1.235686373e-6   ua1 = 2.157228658e-09 lua1 = -6.706068109e-15   ub1 = -1.357459144e-18 lub1 = 1.286205630e-23   uc1 = -3.505848957e-11 luc1 = 5.272007070e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.73 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.114945+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.44751769   k2 = 0.01898311   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.20324992+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7663429+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.0101583   ua = -7.0818604e-10   ub = 1.31832111e-18   uc = -7.1776909e-11   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160310.0   a0 = 1.213479   ags = 0.281809   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -0.0018702   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.14095898   pdiblc1 = 0.39   pdiblc2 = 0.00031929802   pdiblcb = -0.15511953   drout = 0.56   pscbe1 = 799951250.0   pscbe2 = 5.4254628e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.2785893   agidl = 4.4509773e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.88544965   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.4407715   kt2 = -0.052358472   at = 0.0   ute = -0.13226612   ua1 = 1.8227243e-9   ub1 = -7.1588888e-19   uc1 = -8.7612717e-12   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.74 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539359e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584525e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-8   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-07 wpdiblcb = -4.440892099e-22   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 wpscbe2 = 1.323488980e-29 ppscbe2 = 1.058791184e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-7   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23 pub1 = -6.162975822e-45   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.75 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308608e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = -1.387778781e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = 1.110223025e-22 ppclm = -1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343240e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 wuc1 = -1.292469707e-32 puc1 = -2.584939414e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.76 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = -7.112366252e-23 peta0 = -1.387778781e-28   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = -3.330669074e-22 petab = 3.087807787e-28   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493533e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554777e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463398e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16 pagidl = -4.135903063e-37   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = -4.440892099e-22 pute = -2.220446049e-28   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24 pub1 = 6.162975822e-45   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 puc1 = 1.033975766e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.77 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.141052779e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.423581630e-8   k1 = 5.163560651e-01 lk1 = -1.764191989e-10   k2 = -2.646447971e-02 lk2 = 1.698224276e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.340143070e+00 ldsub = -5.902793436e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.023414834e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.817442602e-9   nfactor = {2.915901967e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.323370700e-06 pnfactor = -1.776356839e-27   eta0 = -7.579850000e-02 leta0 = 3.099302733e-7   etab = -1.729996539e+00 letab = 9.473064950e-7   u0 = 1.608035831e-02 lu0 = -6.593709171e-9   ua = 4.365764318e-11 lua = -1.160014925e-15   ub = 1.774933909e-18 lub = 8.121476016e-26   uc = -1.030743287e-10 luc = 4.017669524e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.145642010e+05 lvsat = 1.696810852e-1   a0 = 9.219377220e-01 la0 = -1.125391259e-7   ags = 1.120744390e-01 lags = 6.233271742e-7   a1 = 0.0   a2 = 1.010836186e+00 la2 = -1.136436256e-8   b0 = 0.0   b1 = 0.0   keta = 1.262339765e-02 lketa = -2.757575910e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.658710871e+00 lpclm = -8.933470478e-7   pdiblc1 = 6.967508558e-02 lpdiblc1 = -3.214058779e-8   pdiblc2 = 8.571161110e-04 lpdiblc2 = -4.475215832e-10   pdiblcb = -3.099359191e-02 lpdiblcb = 6.279935762e-9   drout = 1.0   pscbe1 = 7.712957009e+08 lpscbe1 = 1.572349742e+1   pscbe2 = 9.010895465e-09 lpscbe2 = 1.737841029e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.481371233e+00 lbeta0 = 1.243560211e-6   agidl = 8.536887886e-10 lagidl = -3.621444101e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.144215274e-01 lkt1 = -6.773154207e-8   kt2 = -6.597205099e-02 lkt2 = 1.824476986e-8   at = 9.098087549e+04 lat = -3.061507655e-2   ute = -1.978949816e+00 lute = 9.752585094e-7   ua1 = -3.713662156e-09 lua1 = 3.440115825e-15 wua1 = -1.654361225e-30   ub1 = 4.546885644e-18 lub1 = -3.826474399e-24 wub1 = 3.081487911e-39 pub1 = -1.540743956e-45   uc1 = 3.542254351e-10 luc1 = -3.010327285e-16 wuc1 = -2.067951531e-31 puc1 = -2.067951531e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.78 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.074350799e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.301860543e-9   k1 = 4.918287993e-01 lk1 = 1.325900381e-8   k2 = 2.165076081e-02 lk2 = -9.374083109e-09 wk2 = 1.387778781e-23 pk2 = -3.469446952e-30   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -3.943573436e-01 ldsub = 3.598366204e-07 pdsub = 2.220446049e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.975627001e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.002553889e-10   nfactor = {-1.648674244e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.176990034e-06 pnfactor = -4.440892099e-28   eta0 = 0.49   etab = -1.361993125e-03 letab = 4.037064090e-10   u0 = 2.185793948e-03 lu0 = 1.017385823e-9   ua = -3.659750026e-09 lua = 8.686192116e-16   ub = 3.645115856e-18 lub = -9.432241560e-25   uc = -6.519611348e-11 luc = 1.942795591e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.597802425e+05 lvsat = -9.015294234e-2   a0 = 8.634598290e-01 la0 = -8.050639808e-8   ags = 9.193506400e-01 lags = 1.811214532e-7   a1 = 0.0   a2 = 1.216505717e+00 la2 = -1.240249899e-7   b0 = 0.0   b1 = 0.0   keta = -4.296598660e-02 lketa = 2.874715860e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.996019656e-01 lpclm = 3.984777661e-07 wpclm = -3.330669074e-22 ppclm = -1.387778781e-28   pdiblc1 = -4.628132577e-01 lpdiblc1 = 2.595432144e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = -2.081668171e-28   pdiblc2 = -1.086232749e-02 lpdiblc2 = 5.972096636e-09 wpdiblc2 = -5.529431080e-24 ppdiblc2 = 7.318364664e-31   pdiblcb = 2.150677307e-01 lpdiblcb = -1.285063052e-07 wpdiblcb = -5.551115123e-23 ppdiblcb = -1.387778781e-29   drout = 1.608574059e+00 ldrout = -3.333616552e-7   pscbe1 = 8.000344823e+08 lpscbe1 = -1.888856653e-2   pscbe2 = 9.534523798e-09 lpscbe2 = -1.130464069e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.507272163e+00 lbeta0 = 1.338223295e-7   agidl = 3.028298641e-10 lagidl = -6.039766277e-17 wagidl = 4.135903063e-31   bgidl = 6.898757943e+08 lbgidl = 1.698782868e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.626832716e-01 lkt1 = 1.348253482e-8   kt2 = -8.463546509e-03 lkt2 = -1.325695119e-8   at = -8.939633778e+03 lat = 2.411888042e-2   ute = 5.942098076e-01 lute = -4.342540036e-07 pute = 2.220446049e-28   ua1 = 5.277541258e-09 lua1 = -1.485040625e-15   ub1 = -5.135986154e-18 lub1 = 1.477560701e-24   uc1 = -3.045291189e-10 luc1 = 5.981654738e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.79 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.170981582e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.647237095e-8   k1 = -7.903448228e-01 lk1 = 3.950582541e-7   k2 = 4.591602575e-01 lk2 = -1.396534735e-07 wk2 = 5.551115123e-23 pk2 = 9.714451465e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.090266059e-01 ldsub = 1.801639649e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.953485947e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.459560631e-9   nfactor = {4.640460629e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.957571028e-7   eta0 = 7.577509117e-01 leta0 = -7.972952773e-8   etab = -6.25e-6   u0 = 1.677517422e-02 lu0 = -3.326966888e-9   ua = 4.748111728e-09 lua = -1.635031822e-15 wua = -3.308722450e-30   ub = -4.520734203e-18 lub = 1.488361845e-24   uc = 3.218979895e-11 luc = -9.571134166e-18 wuc = -2.039678757e-32 puc = -3.584583953e-39   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -2.156314368e+05 lvsat = 8.119027046e-02 pvsat = -5.820766091e-23   a0 = -4.562594250e-01 la0 = 3.124730028e-7   ags = 2.430890571e+00 lags = -2.689773499e-7   a1 = 0.0   a2 = 1.549941053e+00 la2 = -2.233136970e-7   b0 = 0.0   b1 = 0.0   keta = 2.391484179e-02 lketa = -1.704072281e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.919889609e-01 lpclm = 4.365177795e-8   pdiblc1 = 4.429612748e-01 lpdiblc1 = -1.017379696e-8   pdiblc2 = 6.769843929e-03 lpdiblc2 = 7.216767912e-10   pdiblcb = -4.860480668e-01 lpdiblcb = 8.026845137e-8   drout = 4.874329590e-01 ldrout = 4.861358645e-10   pscbe1 = 7.998768488e+08 lpscbe1 = 2.805077190e-2   pscbe2 = 1.728337771e-08 lpscbe2 = -2.420461381e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.981773089e+00 lbeta0 = 2.903028160e-7   agidl = -3.056660710e-10 lagidl = 1.207972143e-16   bgidl = 2.107586449e+09 lbgidl = -2.522805034e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.491567409e-01 lkt1 = -2.032282784e-8   kt2 = -8.545314104e-02 lkt2 = 9.668625326e-9   at = 1.399712831e+05 lat = -2.022306787e-2   ute = -2.869904438e+00 lute = 5.972726159e-7   ua1 = 6.021704311e-10 lua1 = -9.283207720e-17   ub1 = -1.938790441e-18 lub1 = 5.255157473e-25 pub1 = 1.925929944e-46   uc1 = -3.265376634e-10 luc1 = 6.637014171e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.80 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.12e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-9.391076394e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.830880657e-08 wvth0 = 1.042218585e-12 pvth0 = -2.551090557e-19   k1 = -1.481292926e-02 lk1 = 2.347126300e-07 wk1 = 5.469366471e-13 pk1 = -1.338764175e-19   k2 = 2.758685222e-01 lk2 = -1.052112839e-07 wk2 = 1.442940825e-13 pk2 = -3.531958370e-20   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 5.993096044e+00 ldsub = -1.222185084e-06 wdsub = -7.103845547e-13 pdsub = 1.738843771e-19   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {1.053646952e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.517559055e-08 wvoff = -9.768696785e-14 pvoff = 2.391132758e-20   nfactor = {1.356394467e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.617232141e-08 wnfactor = 2.803651213e-11 pnfactor = -6.862637257e-18   eta0 = 1.881252420e+00 leta0 = -3.606852272e-07 weta0 = -1.086611136e-11 peta0 = 2.659752408e-18   etab = 8.278219153e-02 letab = -2.026454077e-08 wetab = 1.244019324e-12 petab = -3.045048300e-19   u0 = -6.395945592e-03 lu0 = 2.096435602e-09 wu0 = 1.847492978e-14 pu0 = -4.522200940e-21   ua = -5.318116610e-09 lua = 7.068985266e-16 wua = 6.330050830e-21 pua = -1.549438189e-27   ub = 4.052462729e-18 lub = -4.990584633e-25 wub = 2.254913469e-29 pub = -5.519464449e-36   uc = -8.032443944e-11 luc = 1.725519640e-17 wuc = 3.635552862e-22 puc = -8.898924520e-29   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.037548602e+05 lvsat = -1.133153700e-01 wvsat = -7.512069494e-07 pvsat = 1.838766814e-13   a0 = 9.068423576e-01 la0 = 2.141204168e-09 wa0 = 1.260080631e-11 pa0 = -3.084362366e-18   ags = 1.25   a1 = 0.0   a2 = -1.127056235e+00 la2 = 4.152812838e-07 wa2 = -3.168963111e-12 pa2 = 7.756829454e-19   b0 = 0.0   b1 = 0.0   keta = -4.115646522e-01 lketa = 8.828193502e-08 wketa = 1.126831749e-11 pketa = -2.758202413e-18   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.123248131e+00 lpclm = -1.076067325e-07 wpclm = 1.653687455e-12 ppclm = -4.047813480e-19   pdiblc1 = 2.153585552e+00 lpdiblc1 = -4.296511764e-07 wpdiblc1 = -1.574194912e-11 ppdiblc1 = 3.853235596e-18   pdiblc2 = 6.079524328e-02 lpdiblc2 = -1.244852795e-08 wpdiblc2 = 2.302865162e-13 ppdiblc2 = -5.636838199e-20   pdiblcb = 1.325729014e+00 lpdiblcb = -3.572184433e-07 wpdiblcb = 4.894296553e-11 ppdiblcb = -1.198001439e-17   drout = -3.164756316e+00 ldrout = 8.944870484e-07 wdrout = 4.714377852e-11 pdrout = -1.153961839e-17   pscbe1 = 800000000.0   pscbe2 = -5.376496269e-09 lpscbe2 = 2.945458000e-15 wpscbe2 = -2.385549697e-19 ppscbe2 = 5.839229272e-26   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.660750165e+01 lbeta0 = -1.799393126e-06 wbeta0 = 2.871972004e-11 pbeta0 = -7.029869465e-18   agidl = -2.007284338e-09 lagidl = 5.463265326e-16 wagidl = 4.019552251e-19 pagidl = -9.838859023e-26   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.387120560e-01 lkt1 = -4.887372100e-08 wkt1 = 1.136880350e-12 pkt1 = -2.782798880e-19   kt2 = 3.382471888e-01 lkt2 = -9.332100452e-08 wkt2 = 1.940671239e-12 pkt2 = -4.750278024e-19   at = 2.582799737e+05 lat = -5.069142742e-02 wat = -7.111350098e-07 pat = 1.740680720e-13   ute = -1.985225023e+00 lute = 4.253026874e-07 wute = -4.425981796e-12 pute = 1.083369694e-18   ua1 = -3.735522051e-09 lua1 = 9.619980728e-16 wua1 = -3.339909468e-20 pua1 = 8.175263397e-27   ub1 = 6.389055051e-18 lub1 = -1.473710736e-24 wub1 = 3.832196285e-29 pub1 = -9.380258457e-36   uc1 = -1.297570938e-10 luc1 = 2.315671706e-17 wuc1 = 2.682731967e-21 puc1 = -6.566657174e-28   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.81 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.136520303e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.325368137e-7   k1 = 4.276806174e-01 lk1 = 3.976891689e-7   k2 = 4.689033131e-02 lk2 = -5.594776937e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -2.099956519e-06 lcit = 2.425772058e-10 wcit = -1.694065895e-27 pcit = -1.626303259e-31   voff = {-1.783160135e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.998693471e-7   nfactor = {1.703775898e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.254329181e-6   eta0 = 0.08   etab = -0.07   u0 = 7.285540695e-03 lu0 = 5.759243218e-8   ua = -7.222091363e-10 lua = 2.811318801e-16   ub = 4.302881048e-19 lub = 1.780308588e-23 pub = 2.465190329e-44   uc = -1.141547466e-10 luc = 8.495813531e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.006963303e+04 lvsat = 2.009596323e+0   a0 = 1.526779858e+00 la0 = -6.280985109e-6   ags = 7.105961256e-02 lags = 4.225056301e-6   a1 = 0.0   a2 = 1.012601522e+00 la2 = -4.262187475e-6   b0 = 3.429387608e-08 lb0 = -6.875159114e-13   b1 = -5.001763451e-09 lb1 = 1.002742283e-13   keta = 2.968419166e-02 lketa = -6.325953443e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.656496613e-02 lpclm = 3.158004629e-06 ppclm = 1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 1.517196017e-03 lpdiblc2 = -2.401518953e-8   pdiblcb = -2.425118492e-01 lpdiblcb = 1.752021553e-6   drout = 0.56   pscbe1 = 8.000122166e+08 lpscbe1 = -1.222244938e+0   pscbe2 = 1.122218361e-08 lpscbe2 = -1.162113546e-13   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -2.505971875e-11 lalpha0 = 2.507169103e-15   alpha1 = -2.505971875e-11 lalpha1 = 2.507169103e-15   beta0 = 3.594451880e+01 lbeta0 = -5.947358799e-4   agidl = 2.264916321e-09 lagidl = -3.648331365e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = -9.683147321e-02 legidl = 1.969255094e-05 pegidl = 2.131628207e-26   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.376181192e-01 lkt1 = -6.321826893e-8   kt2 = -6.009657711e-02 lkt2 = 1.551317903e-7   at = 8.877989434e+04 lat = -1.779839346e+0   ute = -7.062903695e-02 lute = -1.235686373e-6   ua1 = 2.157228658e-09 lua1 = -6.706068109e-15   ub1 = -1.357459144e-18 lub1 = 1.286205630e-23   uc1 = -3.505848957e-11 luc1 = 5.272007070e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.82 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.114945+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.44751769   k2 = 0.01898311   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.20324992+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7663429+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.0101583   ua = -7.0818604e-10   ub = 1.31832111e-18   uc = -7.1776909e-11   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 160310.0   a0 = 1.213479   ags = 0.281809   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -0.0018702   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.14095898   pdiblc1 = 0.39   pdiblc2 = 0.00031929802   pdiblcb = -0.15511953   drout = 0.56   pscbe1 = 799951250.0   pscbe2 = 5.4254628e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.2785893   agidl = 4.4509773e-10   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.88544965   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.4407715   kt2 = -0.052358472   at = 0.0   ute = -0.13226612   ua1 = 1.8227243e-9   ub1 = -7.1588888e-19   uc1 = -8.7612717e-12   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.83 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539359e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584524e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-8   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 ppscbe2 = 2.117582368e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-07 wute = 4.440892099e-22   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23 pub1 = -1.232595164e-44   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.84 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308608e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = -2.775557562e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = 2.220446049e-22 ppclm = -4.440892099e-28   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14 wpscbe2 = -1.058791184e-28   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343240e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 puc1 = 5.169878828e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.85 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-06 pdsub = -8.881784197e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = 8.673617380e-23 peta0 = -4.007211230e-28   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = 6.990935608e-22 petab = -1.377370440e-27   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493533e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554777e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463397e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-07 wpdiblc1 = 1.776356839e-21   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16 pagidl = 8.271806126e-37   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = 4.440892099e-22 pute = -4.440892099e-28   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24 pub1 = -6.162975822e-45   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 puc1 = -1.033975766e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.86 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.141052779e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.423581630e-8   k1 = 5.163560651e-01 lk1 = -1.764191989e-10   k2 = -2.646447971e-02 lk2 = 1.698224276e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.340143070e+00 ldsub = -5.902793436e-07 pdsub = 1.776356839e-27   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.023414834e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.817442602e-9   nfactor = {2.915901967e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.323370700e-06 wnfactor = 7.105427358e-21   eta0 = -7.579850000e-02 leta0 = 3.099302733e-7   etab = -1.729996539e+00 letab = 9.473064950e-7   u0 = 1.608035831e-02 lu0 = -6.593709171e-9   ua = 4.365764318e-11 lua = -1.160014925e-15   ub = 1.774933909e-18 lub = 8.121476016e-26   uc = -1.030743287e-10 luc = 4.017669524e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.145642010e+05 lvsat = 1.696810852e-1   a0 = 9.219377220e-01 la0 = -1.125391259e-7   ags = 1.120744390e-01 lags = 6.233271742e-7   a1 = 0.0   a2 = 1.010836186e+00 la2 = -1.136436256e-8   b0 = 0.0   b1 = 0.0   keta = 1.262339765e-02 lketa = -2.757575910e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.658710871e+00 lpclm = -8.933470478e-7   pdiblc1 = 6.967508558e-02 lpdiblc1 = -3.214058779e-8   pdiblc2 = 8.571161110e-04 lpdiblc2 = -4.475215832e-10   pdiblcb = -3.099359191e-02 lpdiblcb = 6.279935762e-9   drout = 1.0   pscbe1 = 7.712957009e+08 lpscbe1 = 1.572349742e+1   pscbe2 = 9.010895465e-09 lpscbe2 = 1.737841029e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.481371233e+00 lbeta0 = 1.243560211e-6   agidl = 8.536887886e-10 lagidl = -3.621444101e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.144215274e-01 lkt1 = -6.773154207e-8   kt2 = -6.597205099e-02 lkt2 = 1.824476986e-8   at = 9.098087549e+04 lat = -3.061507655e-2   ute = -1.978949816e+00 lute = 9.752585094e-7   ua1 = -3.713662156e-09 lua1 = 3.440115825e-15 wua1 = -1.654361225e-30 pua1 = -2.481541838e-36   ub1 = 4.546885644e-18 lub1 = -3.826474399e-24 wub1 = 6.162975822e-39 pub1 = -3.081487911e-45   uc1 = 3.542254351e-10 luc1 = -3.010327285e-16 puc1 = -2.067951531e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.87 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.074350799e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.301860543e-9   k1 = 4.918287993e-01 lk1 = 1.325900381e-8   k2 = 2.165076081e-02 lk2 = -9.374083109e-09 pk2 = 1.387778781e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -3.943573436e-01 ldsub = 3.598366204e-07 pdsub = 4.440892099e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.975627001e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.002553889e-10   nfactor = {-1.648674244e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.176990034e-06 pnfactor = -8.881784197e-28   eta0 = 0.49   etab = -1.361993125e-03 letab = 4.037064090e-10   u0 = 2.185793948e-03 lu0 = 1.017385823e-9   ua = -3.659750026e-09 lua = 8.686192116e-16   ub = 3.645115856e-18 lub = -9.432241560e-25   uc = -6.519611348e-11 luc = 1.942795591e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.597802425e+05 lvsat = -9.015294234e-2   a0 = 8.634598290e-01 la0 = -8.050639808e-8   ags = 9.193506400e-01 lags = 1.811214532e-7   a1 = 0.0   a2 = 1.216505717e+00 la2 = -1.240249899e-07 wa2 = 3.552713679e-21   b0 = 0.0   b1 = 0.0   keta = -4.296598660e-02 lketa = 2.874715860e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.996019656e-01 lpclm = 3.984777661e-07 wpclm = -1.110223025e-22 ppclm = 8.326672685e-29   pdiblc1 = -4.628132577e-01 lpdiblc1 = 2.595432144e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = -2.220446049e-28   pdiblc2 = -1.086232749e-02 lpdiblc2 = 5.972096636e-09 wpdiblc2 = -1.235990477e-23 ppdiblc2 = -8.673617380e-31   pdiblcb = 2.150677307e-01 lpdiblcb = -1.285063052e-07 wpdiblcb = -1.110223025e-22 ppdiblcb = -1.110223025e-28   drout = 1.608574059e+00 ldrout = -3.333616552e-7   pscbe1 = 8.000344823e+08 lpscbe1 = -1.888856653e-2   pscbe2 = 9.534523798e-09 lpscbe2 = -1.130464069e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.507272163e+00 lbeta0 = 1.338223295e-7   agidl = 3.028298641e-10 lagidl = -6.039766277e-17   bgidl = 6.898757943e+08 lbgidl = 1.698782868e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.626832716e-01 lkt1 = 1.348253482e-8   kt2 = -8.463546509e-03 lkt2 = -1.325695119e-8   at = -8.939633778e+03 lat = 2.411888042e-2   ute = 5.942098076e-01 lute = -4.342540036e-07 pute = -2.220446049e-28   ua1 = 5.277541258e-09 lua1 = -1.485040625e-15 pua1 = 3.308722450e-36   ub1 = -5.135986154e-18 lub1 = 1.477560701e-24   uc1 = -3.045291189e-10 luc1 = 5.981654738e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.25e-6   sbref = 1.24e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.88 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.170981583e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.647237095e-8   k1 = -7.903448228e-01 lk1 = 3.950582541e-7   k2 = 4.591602575e-01 lk2 = -1.396534735e-07 wk2 = 1.110223025e-22 pk2 = 8.326672685e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.090266059e-01 ldsub = 1.801639649e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.953485947e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.459560631e-9   nfactor = {4.640460629e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.957571028e-7   eta0 = 7.577509117e-01 leta0 = -7.972952773e-8   etab = -6.25e-6   u0 = 1.677517422e-02 lu0 = -3.326966888e-9   ua = 4.748111728e-09 lua = -1.635031822e-15 wua = -6.617444900e-30   ub = -4.520734203e-18 lub = 1.488361845e-24 wub = 6.162975822e-39 pub = -7.703719778e-46   uc = 3.218979895e-11 luc = -9.571134166e-18 wuc = 3.635071051e-33 puc = -1.090521315e-38   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -2.156314368e+05 lvsat = 8.119027046e-02 pvsat = -1.164153218e-22   a0 = -4.562594250e-01 la0 = 3.124730028e-7   ags = 2.430890571e+00 lags = -2.689773499e-7   a1 = 0.0   a2 = 1.549941053e+00 la2 = -2.233136970e-7   b0 = 0.0   b1 = 0.0   keta = 2.391484179e-02 lketa = -1.704072281e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.919889609e-01 lpclm = 4.365177795e-8   pdiblc1 = 4.429612748e-01 lpdiblc1 = -1.017379696e-8   pdiblc2 = 6.769843929e-03 lpdiblc2 = 7.216767912e-10   pdiblcb = -4.860480668e-01 lpdiblcb = 8.026845137e-8   drout = 4.874329590e-01 ldrout = 4.861358645e-10   pscbe1 = 7.998768488e+08 lpscbe1 = 2.805077190e-2   pscbe2 = 1.728337771e-08 lpscbe2 = -2.420461381e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.981773089e+00 lbeta0 = 2.903028160e-7   agidl = -3.056660710e-10 lagidl = 1.207972143e-16   bgidl = 2.107586449e+09 lbgidl = -2.522805034e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.491567409e-01 lkt1 = -2.032282784e-8   kt2 = -8.545314104e-02 lkt2 = 9.668625326e-9   at = 1.399712831e+05 lat = -2.022306787e-2   ute = -2.869904438e+00 lute = 5.972726159e-07 pute = 1.776356839e-27   ua1 = 6.021704311e-10 lua1 = -9.283207720e-17   ub1 = -1.938790441e-18 lub1 = 5.255157473e-25 pub1 = 3.851859889e-46   uc1 = -3.265376634e-10 luc1 = 6.637014171e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.89 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 9.4e-07 wmax = 1.0e-6   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-8.746854723e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.367687654e-07 wvth0 = -7.973307283e-07 pvth0 = 1.951666290e-13   k1 = 1.128011385e+00 lk1 = -4.502219149e-08 wk1 = -1.069948146e-06 pk1 = 2.618965575e-13   k2 = -1.621327355e+00 lk2 = 3.591748369e-07 wk2 = 1.776215634e-06 pk2 = -4.347731819e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 6.244505849e+00 ldsub = -1.283723919e-06 wdsub = -2.353786145e-07 pdsub = 5.761480036e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {6.912619995e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.185886032e-07 wvoff = -5.485359027e-07 pvoff = 1.342678756e-13   nfactor = {1.635226799e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.614442620e-06 wnfactor = -1.403958862e-05 pnfactor = 3.436540305e-12   eta0 = 2.492190326e+00 leta0 = -5.102275532e-07 weta0 = -5.719904838e-07 peta0 = 1.400089707e-13   etab = -4.693748349e-01 letab = 1.148896954e-07 wetab = 5.169483212e-07 petab = -1.265360253e-13   u0 = 2.135825079e-02 lu0 = -4.697097816e-09 wu0 = -2.598434831e-08 pu0 = 6.360318857e-15   ua = 3.347872427e-08 lua = -8.789598200e-15 wua = -3.632283760e-14 pua = 8.890922574e-21   ub = -3.370901887e-17 lub = 8.744008196e-24 wub = 3.535352999e-23 pub = -8.653660304e-30   uc = -7.789411672e-11 luc = 1.666031415e-17 wuc = -2.274982350e-18 puc = 5.568588048e-25   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.324122118e+07 lvsat = -1.299765119e+01 wvsat = -4.928088112e+01 pvsat = 1.206272768e-5   a0 = 8.426059942e+00 la0 = -1.838375280e-06 wa0 = -7.039719517e-06 pa0 = 1.723147345e-12   ags = 1.250000033e+00 lags = -8.198270507e-15 wags = -3.135730253e-14 pags = 7.675478031e-21   a1 = 0.0   a2 = -6.764742225e+00 la2 = 1.795245872e-06 wa2 = 5.278178860e-06 pa2 = -1.291966230e-12   b0 = 0.0   b1 = 0.0   keta = -3.665176758e-01 lketa = 7.725556137e-08 wketa = -4.216315249e-08 pketa = 1.032048565e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.117998897e+00 lpclm = -1.063218512e-07 wpclm = 4.916154842e-09 ppclm = -1.203351801e-15   pdiblc1 = 2.664329522e+00 lpdiblc1 = -5.546685315e-07 wpdiblc1 = -4.781905897e-07 ppdiblc1 = 1.170491016e-13   pdiblc2 = 9.660757903e-02 lpdiblc2 = -2.121449243e-08 wpdiblc2 = -3.352842443e-08 ppdiblc2 = 8.206920091e-15   pdiblcb = -1.487182724e-01 lpdiblcb = 3.689391366e-09 wpdiblcb = 1.380473675e-06 ppdiblcb = -3.379054439e-13   drout = -3.164706465e+00 ldrout = 8.944748462e-07 wdrout = 4.722523528e-13 pdrout = -1.155955687e-19   pscbe1 = 7.999999948e+08 lpscbe1 = 1.266220093e-06 wpscbe1 = 4.843139648e-06 ppscbe1 = -1.185478210e-12   pscbe2 = -3.891186874e-08 lpscbe2 = 1.115407880e-14 wpscbe2 = 3.139665029e-14 ppscbe2 = -7.685115074e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 2.087149899e+01 lbeta0 = -2.843113073e-06 wbeta0 = -3.992062032e-06 pbeta0 = 9.771569839e-13   agidl = -5.801812013e-08 lagidl = 1.425637886e-14 wagidl = 5.243953877e-14 pagidl = -1.283588810e-20   bgidl = 9.999999963e+08 lbgidl = 9.019279480e-07 wbgidl = 3.449752808e-06 pbgidl = -8.444099426e-13   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 7.032593021e-01 lkt1 = -3.039222602e-07 wkt1 = -9.755257916e-07 pkt1 = 2.387843256e-13   kt2 = 3.382492550e-01 lkt2 = -9.332151027e-08 wkt2 = 6.217426574e-15 pkt2 = -1.521870185e-21   at = 9.223499639e+05 lat = -2.132391593e-01 wat = -6.217242861e-01 pat = 1.521825621e-7   ute = -3.558028776e+00 lute = 8.102857261e-07 wute = 1.472504778e-06 pute = -3.604323570e-13   ua1 = -3.735557882e-09 lua1 = 9.620068433e-16 wua1 = 1.470091689e-22 pua1 = -3.598416983e-29   ub1 = 6.389096846e-18 lub1 = -1.473720966e-24 wub1 = -8.076284485e-31 pub1 = 1.976872517e-37   uc1 = -1.297542173e-10 luc1 = 2.315601297e-17 wuc1 = -1.032124205e-23 puc1 = 2.526382058e-30   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.90 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.179549702e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.737532466e-06 wvth0 = 3.770373655e-08 pvth0 = -3.772174951e-12   k1 = 3.881179132e-01 lk1 = 4.355849698e-06 wk1 = 3.466610743e-08 pk1 = -3.468266916e-12   k2 = 1.025479962e-01 lk2 = -6.127903231e-06 wk2 = -4.876902705e-08 pk2 = 4.879232645e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -2.623189420e-05 lcit = 2.656923877e-09 wcit = 2.114517602e-11 pcit = -2.115527813e-15   voff = {-1.285882747e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.475018972e-06 wvoff = -4.357303604e-08 pvoff = 4.359385306e-12   nfactor = {1.578993384e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.373854208e-05 wnfactor = 1.093384320e-07 pnfactor = -1.093906684e-11   eta0 = 0.08   etab = -0.07   u0 = 1.556160723e-03 lu0 = 6.308041505e-07 wu0 = 5.020266071e-09 pu0 = -5.022664503e-13   ua = -7.501765498e-10 lua = 3.079209370e-15 wua = 2.450594264e-17 pua = -2.451765035e-21   ub = -1.340789098e-18 lub = 1.949954193e-22 wub = 1.551874519e-24 pub = -1.552615927e-28   uc = -1.986723508e-10 luc = 9.305379602e-15 wuc = 7.405702937e-17 puc = -7.409241011e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.398479688e+05 lvsat = 2.201090756e+01 wvsat = 1.751742000e-01 pvsat = -1.752578895e-5   a0 = 2.151621507e+00 la0 = -6.879500180e-05 wa0 = -5.475062476e-07 pa0 = 5.477678187e-11   ags = -3.492552106e-01 lags = 4.627661916e-05 wags = 3.682932981e-07 pags = -3.684692502e-11   a1 = 0.0   a2 = 1.436610209e+00 la2 = -4.668331320e-05 wa2 = -3.715299799e-07 pa2 = 3.717074783e-11   b0 = 1.026889715e-07 lb0 = -7.530293026e-12 wb0 = -5.992997123e-14 pb0 = 5.995860277e-18   b1 = -1.497719136e-08 lb1 = 1.098293595e-12 wb1 = 8.740789144e-15 pb1 = -8.744965057e-19   keta = 9.261570815e-02 lketa = -6.928753547e-06 wketa = -5.514260856e-08 pketa = 5.516895294e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -3.307279175e-01 lpclm = 3.458930890e-05 wpclm = 2.752796312e-07 ppclm = -2.754111461e-11   pdiblc1 = 0.39   pdiblc2 = 3.906262439e-03 lpdiblc2 = -2.630359694e-07 wpdiblc2 = -2.093376449e-09 ppdiblc2 = 2.094376560e-13   pdiblcb = -4.168055336e-01 lpdiblcb = 1.918971687e-05 wpdiblcb = 1.527217036e-07 ppdiblcb = -1.527946664e-11   drout = 0.56   pscbe1 = 8.001338073e+08 lpscbe1 = -1.338712658e+01 wpscbe1 = -1.065416854e-01 ppscbe1 = 1.065925857e-5   pscbe2 = 2.278306031e-08 lpscbe2 = -1.272851345e-12 wpscbe2 = -1.013001011e-14 ppscbe2 = 1.013484972e-18   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -2.744765935e-10 lalpha0 = 2.746077247e-14 walpha0 = 2.185470470e-16 palpha0 = -2.186514578e-20   alpha1 = -2.744765935e-10 lalpha1 = 2.746077247e-14 walpha1 = 2.185470470e-16 palpha1 = -2.186514578e-20   beta0 = 9.510972002e+01 lbeta0 = -6.514082619e-03 wbeta0 = -5.184244259e-05 pbeta0 = 5.186721032e-9   agidl = 5.894330092e-09 lagidl = -3.995980860e-13 wagidl = -3.180208488e-15 pagidl = 3.181727832e-19   bgidl = 1000000000.0   cgidl = 300.0   egidl = -2.055875443e+00 legidl = 2.156905412e-04 wegidl = 1.716577016e-06 pegidl = -1.717397110e-10   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.313290727e-01 lkt1 = -6.924233778e-07 wkt1 = -5.510663790e-09 pkt1 = 5.513296510e-13   kt2 = -7.552931608e-02 lkt2 = 1.699142986e-06 wkt2 = 1.352265973e-08 pkt2 = -1.352912018e-12   at = 2.658409337e+05 lat = -1.949440238e+01 wat = -1.551465487e-01 pat = 1.552206699e-5   ute = 5.229886324e-02 lute = -1.353434927e-05 wute = -1.077133598e-07 pute = 1.077648199e-11   ua1 = 2.824358190e-09 lua1 = -7.345089339e-14 wua1 = -5.845602438e-16 pua1 = 5.848395174e-20   ub1 = -2.636995446e-18 lub1 = 1.408768164e-22 wub1 = 1.121170654e-24 pub1 = -1.121706293e-28   uc1 = -8.750519233e-11 luc1 = 5.774376624e-15 wuc1 = 4.595547925e-17 puc1 = -4.597743448e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.91 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-8.280823385e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.308606156e-06 wvth0 = -2.513582436e-07 pvth0 = 2.022874589e-12   k1 = 7.112690514e-01 lk1 = -2.122611612e-06 wk1 = -2.311073829e-07 pk1 = 1.859900218e-12   k2 = -3.520679895e-01 lk2 = 2.986135762e-06 wk2 = 3.251268470e-07 pk2 = -2.616547711e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.708795846e-04 lcit = -1.294722699e-09 wcit = -1.409678401e-10 pcit = 1.134477460e-15   voff = {-5.347681788e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.667984355e-06 wvoff = 2.904869069e-07 pvoff = -2.337773268e-12   nfactor = {2.598226328e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.694810654e-06 wnfactor = -7.289228798e-07 pnfactor = 5.866207329e-12   eta0 = 0.08   etab = -0.07   u0 = 4.835416648e-02 lu0 = -3.073917393e-07 wu0 = -3.346844047e-08 pu0 = 2.693464785e-13   ua = -5.217366169e-10 lua = -1.500503006e-15 wua = -1.633729509e-16 pua = 1.314788750e-21   ub = 1.312550246e-17 lub = -9.502153889e-23 wub = -1.034583013e-23 pub = 8.326091306e-29   uc = 4.916737857e-10 luc = -4.534524415e-15 wuc = -4.937135291e-16 puc = 3.973295397e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.493094012e+06 lvsat = -1.072594585e+01 wvsat = -1.167828000e+00 pvsat = 9.398416985e-6   a0 = -2.952131992e+00 la0 = 3.352390000e-05 wa0 = 3.650041651e-06 pa0 = -2.937471395e-11   ags = 3.083907821e+00 lags = -2.255066084e-05 wags = -2.455288654e-06 pags = 1.975961065e-11   a1 = 0.0   a2 = -2.026724580e+00 la2 = 2.274884341e-05 wa2 = 2.476866533e-06 pa2 = -1.993326456e-11   b0 = -4.559673026e-07 lb0 = 3.669522259e-12 wb0 = 3.995331415e-13 pb0 = -3.215352828e-18   b1 = 6.650285270e-08 lb1 = -5.351999954e-13 wb1 = -5.827192763e-14 pb1 = 4.689593624e-19   keta = -4.214136433e-01 lketa = 3.376391234e-06 wketa = 3.676173904e-07 pketa = -2.958502044e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.235378656e+00 lpclm = -1.685541831e-05 wpclm = -1.835197541e-06 ppclm = 1.476925689e-11   pdiblc1 = 0.39   pdiblc2 = -1.560781146e-02 lpdiblc2 = 1.281777935e-07 wpdiblc2 = 1.395584299e-08 ppdiblc2 = -1.123134843e-13   pdiblcb = 1.006838366e+00 lpdiblcb = -9.351175703e-06 wpdiblcb = -1.018144691e-06 ppdiblcb = 8.193799388e-12   drout = 0.56   pscbe1 = 7.991406452e+08 lpscbe1 = 6.523565390e+00 wpscbe1 = 7.102779027e-01 ppscbe1 = -5.716156749e-6   pscbe2 = -7.164704852e-08 lpscbe2 = 6.202622298e-13 wpscbe2 = 6.753340074e-14 ppscbe2 = -5.434936142e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.762779165e-09 lalpha0 = -1.338167259e-14 walpha0 = -1.456980313e-15 palpha0 = 1.172544974e-20   alpha1 = 1.762779165e-09 lalpha1 = -1.338167259e-14 walpha1 = -1.456980313e-15 palpha1 = 1.172544974e-20   beta0 = -3.881560855e+02 lbeta0 = 3.174321515e-03 wbeta0 = 3.456162839e-04 pbeta0 = -2.781442089e-9   agidl = -2.375099408e-08 lagidl = 1.947247028e-13 wagidl = 2.120138992e-14 pagidl = -1.706240158e-19   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.394574278e+01 legidl = -1.051063006e-04 wegidl = -1.144384677e-05 pegidl = 9.209750395e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.826984766e-01 lkt1 = 3.374188745e-07 wkt1 = 3.673775860e-08 pkt1 = -2.956572152e-13   kt2 = 5.052645441e-02 lkt2 = -8.279947386e-07 wkt2 = -9.015106484e-08 pkt2 = 7.255154858e-13   at = -1.180406929e+06 lat = 9.499649375e+00 wat = 1.034310324e+00 pat = -8.323896771e-6   ute = -9.517854546e-01 lute = 6.595307213e-06 wute = 7.180890656e-07 pute = -5.779019230e-12   ua1 = -2.624805911e-09 lua1 = 3.579272244e-14 wua1 = 3.897068292e-15 pua1 = -3.136272877e-20   ub1 = 7.814353137e-18 lub1 = -6.864946845e-23 wub1 = -7.474471023e-24 pub1 = 6.015286104e-29   uc1 = 3.408834133e-10 luc1 = -2.813861755e-15 wuc1 = -3.063698617e-16 puc1 = 2.465595713e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.92 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539359e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584524e+05 lvsat = -8.703544119e-01 wvsat = 4.656612873e-16   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-8   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 ppscbe2 = 5.293955920e-35   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-7   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.93 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308607e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = 1.387778781e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = 2.220446049e-22 ppclm = -1.110223025e-27   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343240e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 puc1 = 2.584939414e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.94 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-06 pdsub = -8.881784197e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = -6.938893904e-23 peta0 = 1.040834086e-29   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = -5.204170428e-24 petab = 5.967448757e-28   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493534e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554778e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463398e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16 pagidl = -4.135903063e-37   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = -8.881784197e-22 pute = 8.881784197e-28   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15 pua1 = 6.617444900e-36   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24 pub1 = -6.162975822e-45   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 puc1 = -1.033975766e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.95 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.150304223e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.392924790e-08 wvth0 = 8.106411162e-09 pvth0 = -8.493694956e-15   k1 = 4.478016515e-01 lk1 = 7.165318145e-08 wk1 = 6.006957088e-08 pk1 = -6.293939463e-14   k2 = -1.678314146e-01 lk2 = 1.651029830e-07 wk2 = 1.238702321e-07 pk2 = -1.297881324e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.963615285e+00 ldsub = -1.243537943e-06 wdsub = -5.463063057e-07 pdsub = 5.724060894e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.986018969e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.026766974e-07 wvoff = 8.434645466e-08 pvoff = -8.837610653e-14   nfactor = {2.013559503e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.936573460e-05 wnfactor = -1.508844609e-05 pnfactor = 1.580929660e-11   eta0 = -4.831572070e-01 leta0 = 7.367505426e-07 weta0 = 3.569407345e-07 peta0 = -3.739935781e-13   etab = -1.730313590e+00 letab = 9.476386927e-07 wetab = 2.778099028e-10 petab = -2.910822709e-16   u0 = 3.780880286e-02 lu0 = -2.936023015e-08 wu0 = -1.903915842e-08 pu0 = 1.994875421e-14   ua = 9.567328185e-09 lua = -1.113867883e-14 wua = -8.344944886e-15 pua = 8.743624628e-21   ub = -5.716345550e-18 lub = 7.930390094e-24 wub = 6.564098782e-24 pub = -6.877698601e-30   uc = -1.188024463e-10 luc = 5.665622373e-17 wuc = 1.378148001e-17 puc = -1.443989021e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.265837302e+05 lvsat = 7.061623474e-01 wvsat = 4.486478961e-01 pvsat = -4.700820493e-7   a0 = 1.258262881e+00 la0 = -4.649322190e-07 wa0 = -2.946988664e-07 pa0 = 3.087781047e-13   ags = 1.120744384e-01 lags = 6.233271749e-07 wags = 5.643752132e-16 pags = -5.913403101e-22   a1 = 0.0   a2 = 5.898622379e-01 la2 = 4.297216159e-07 wa2 = 3.688708445e-07 pa2 = -3.864936491e-13   b0 = 9.563527155e-16 lb0 = -1.002042467e-21 wb0 = -8.379868526e-22 pb0 = 8.780216745e-28   b1 = 3.975996046e-19 lb1 = -4.165949258e-25 wb1 = -3.483894968e-25 pb1 = 3.650338050e-31   keta = 7.708845154e-03 lketa = -2.242641386e-08 wketa = 4.306288163e-09 pketa = -4.512021080e-15   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.000827725e+00 lpclm = -1.251808535e-06 wpclm = -2.997737352e-07 ppclm = 3.140954254e-13   pdiblc1 = 1.194479363e-01 lpdiblc1 = -8.429133646e-08 wpdiblc1 = -4.361256454e-08 ppdiblc1 = 4.569615481e-14   pdiblc2 = 1.502606527e-03 lpdiblc2 = -1.123850304e-09 wpdiblc2 = -5.655993580e-10 ppdiblc2 = 5.926208673e-16   pdiblcb = -2.047072165e-01 lpdiblcb = 1.882927288e-07 wpdiblcb = 1.522134367e-07 ppdiblcb = -1.594854337e-13   drout = 5.874033614e-01 ldrout = 4.323084430e-07 wdrout = 3.615303778e-07 pdrout = -3.788024916e-13   pscbe1 = 2.118540502e+08 lpscbe1 = 6.018924730e+02 wpscbe1 = 4.902006765e+02 ppscbe1 = -5.136200139e-4   pscbe2 = 6.721677170e-08 lpscbe2 = -6.081287787e-14 wpscbe2 = -5.100185135e-14 ppscbe2 = 5.343846479e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.219746654e+00 lbeta0 = 1.517683904e-06 wbeta0 = 2.292438281e-07 pbeta0 = -2.401959520e-13   agidl = -1.246073848e-09 lagidl = 1.837934386e-15 wagidl = 1.839879215e-15 pagidl = -1.927779444e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.686070419e-01 lkt1 = -1.157348146e-07 wkt1 = -4.014411822e-08 pkt1 = 4.206200347e-14   kt2 = -8.869667737e-02 lkt2 = 4.205506526e-08 wkt2 = 1.991204482e-08 pkt2 = -2.086334276e-14   at = 1.289488170e+05 lat = -7.039693646e-02 wat = -3.326872532e-02 pat = 3.485813867e-8   ute = -2.012809748e+00 lute = 1.010736099e-06 wute = 2.966915524e-08 pute = -3.108659913e-14   ua1 = -4.475320590e-09 lua1 = 4.238162490e-15 wua1 = 6.673894923e-16 pua1 = -6.992740253e-22   ub1 = 5.876055253e-18 lub1 = -5.219145085e-24 wub1 = -1.164660944e-24 pub1 = 1.220302621e-30   uc1 = 4.624259075e-10 luc1 = -4.144024784e-16 wuc1 = -9.480871633e-17 puc1 = 9.933820275e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.96 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-9.807205760e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.896443411e-08 wvth0 = -8.204179772e-08 pvth0 = 4.088724016e-14   k1 = 1.121012948e+00 lk1 = -2.971151365e-07 wk1 = -5.513112850e-07 pk1 = 2.719597537e-13   k2 = 3.035501063e-02 lk2 = 5.654141388e-08 wk2 = -7.626942235e-09 pk2 = -5.775726776e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -1.990661375e+00 ldsub = 9.225159537e-07 wdsub = 1.398732674e-06 pdsub = -4.930376376e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.588943386e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.218612205e-08 wvoff = -1.591879294e-07 pvoff = 4.502594072e-14   nfactor = {-3.683864771e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.184333122e-05 wnfactor = 3.083458083e-05 pnfactor = -9.346189468e-12   eta0 = 1.304717420e+00 leta0 = -2.426024814e-07 weta0 = -7.138814746e-07 peta0 = 2.125760575e-13   etab = -1.505034174e-03 letab = 6.405860321e-10 wetab = 1.253371447e-10 petab = -2.075615058e-16   u0 = -4.613443752e-02 lu0 = 1.662177834e-08 wu0 = 4.233973306e-08 pu0 = -1.367306807e-14   ua = -2.402105691e-08 lua = 7.260198818e-15 wua = 1.784122865e-14 pua = -5.600506582e-21   ub = 1.976849459e-17 lub = -6.029568213e-24 wub = -1.412782040e-23 pub = 4.456817426e-30   uc = -4.603851097e-11 luc = 1.679795903e-17 wuc = -1.678650437e-17 puc = 2.304487428e-24   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.231791743e+06 lvsat = -8.595842775e-01 wvsat = -1.640316381e+00 pvsat = 6.742003576e-7   a0 = 4.473788908e-01 la0 = -2.075024144e-08 wa0 = 3.645834327e-07 pa0 = -5.236025664e-14   ags = 6.685898265e-01 lags = 3.184819581e-07 wags = 2.197246492e-07 pags = -1.203596700e-13   a1 = 0.0   a2 = 2.011294128e+00 la2 = -3.489032375e-07 wa2 = -6.964190388e-07 pa2 = 1.970455167e-13   b0 = -1.912705431e-15 lb0 = 5.695558597e-22 wb0 = 1.675973705e-21 pb0 = -4.990630701e-28   b1 = -7.951992093e-19 lb1 = 2.367904445e-25 wb1 = 6.967789936e-25 pb1 = -2.074833648e-31   keta = -1.438763007e-02 lketa = -1.032251714e-08 wketa = -2.504127050e-08 pketa = 1.156383786e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.400206340e+00 lpclm = 6.111929001e-07 wpclm = 6.138919719e-07 ppclm = -1.863878073e-13   pdiblc1 = -6.117395955e-01 lpdiblc1 = 3.162349138e-07 wpdiblc1 = 1.304940228e-07 ppdiblc1 = -4.967508107e-14   pdiblc2 = -1.946655045e-02 lpdiblc2 = 1.036252966e-08 wpdiblc2 = 7.539295491e-09 ppdiblc2 = -3.847037909e-15   pdiblcb = -2.855159746e-01 lpdiblcb = 2.325577463e-07 wpdiblcb = 4.386274612e-07 ppdiblcb = -3.163758759e-13   drout = 2.903407127e+00 ldrout = -8.363405196e-07 wdrout = -1.134574169e-06 pdrout = 4.407261763e-13   pscbe1 = 1.918944405e+09 lpscbe1 = -3.332089460e+02 wpscbe1 = -9.804246792e+02 ppscbe1 = 2.919517904e-4   pscbe2 = -1.105542407e-07 lpscbe2 = 3.656563843e-14 wpscbe2 = 1.052256183e-13 ppscbe2 = -3.213903737e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.476501556e+00 lbeta0 = 2.814899877e-07 wbeta0 = 2.696218976e-08 pbeta0 = -1.293911275e-13   agidl = 3.302029760e-09 lagidl = -6.534030676e-16 wagidl = -2.627994923e-15 pagidl = 5.196103119e-22   bgidl = 4.546810828e+08 lbgidl = 2.987120699e+02 wbgidl = 2.060851325e+02 pbgidl = -1.128882834e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -7.168979821e-01 lkt1 = 7.505025515e-08 wkt1 = 1.351278642e-07 pkt1 = -5.394760672e-14   kt2 = 3.900563629e-02 lkt2 = -2.789706960e-08 wkt2 = -4.159401698e-08 pkt2 = 1.282814024e-14   at = -1.343064844e+05 lat = 7.380773629e-02 wat = 1.098504463e-01 pat = -4.353896556e-8   ute = 1.012016512e+00 lute = -6.461881057e-07 wute = -3.660956046e-07 pute = 1.857034422e-13   ua1 = 6.855606336e-09 lua1 = -1.968636007e-15 wua1 = -1.382751119e-15 pua1 = 4.237417483e-22   ub1 = -7.739071597e-18 lub1 = 2.238881025e-24 wub1 = 2.280906763e-24 pub1 = -6.670932301e-31   uc1 = -4.525893734e-10 luc1 = 8.682001708e-17 wuc1 = 1.297351329e-16 puc1 = -2.366130426e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.97 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-2.150135287e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.992580315e-07 wvth0 = 8.579658089e-07 pvth0 = -2.390235249e-13   k1 = 2.848942155e+00 lk1 = -8.116492562e-07 wk1 = -3.188859707e-06 pk1 = 1.057355735e-12   k2 = -1.035043383e+00 lk2 = 3.737904207e-07 wk2 = 1.309269045e-06 pk2 = -4.498959703e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.089764971e+01 ldsub = 6.552544406e-06 wdsub = 1.849434520e-05 pdsub = -5.583683658e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-9.996168260e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.407433022e-07 wvoff = 7.047255609e-07 pvoff = -2.122258989e-13   nfactor = {2.234193947e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.779168130e-06 wnfactor = -1.551060221e-05 pnfactor = 4.454247411e-12   eta0 = -5.338381886e+00 leta0 = 1.735546414e-06 weta0 = 5.341626633e-06 peta0 = -1.590602869e-12   etab = -8.833848892e-01 letab = 2.632423599e-07 wetab = 7.740446318e-07 petab = -2.306613795e-13   u0 = 1.484572263e-01 lu0 = -4.132275436e-08 wu0 = -1.153840279e-07 pu0 = 3.329312485e-14   ua = 5.868115416e-08 lua = -1.736645208e-14 wua = -4.725785763e-14 pua = 1.378437384e-20   ub = -5.302888836e-17 lub = 1.564767249e-23 wub = 4.250439693e-23 pub = -1.240684109e-29   uc = 3.972586092e-10 luc = -1.152048409e-16 wuc = -3.198849737e-16 puc = 9.255963414e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -5.290413727e+06 lvsat = 1.380340456e+00 wvsat = 4.446686635e+00 pvsat = -1.138356966e-6   a0 = 5.678182421e+00 la0 = -1.578352763e-06 wa0 = -5.375194247e-06 pa0 = 1.656802042e-12   ags = 3.326465188e+00 lags = -4.729668775e-07 wags = -7.847311371e-07 pags = 1.787421518e-13   a1 = 0.0   a2 = 4.169311456e+00 la2 = -9.915068476e-07 wa2 = -2.295176168e-06 pa2 = 6.731154207e-13   b0 = 0.0   b1 = 0.0   keta = 1.630440660e+00 lketa = -5.001112612e-07 wketa = -1.407689331e-06 pketa = 4.232818640e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.443110656e+00 lpclm = 6.239687330e-07 wpclm = 1.695596208e-06 ppclm = -5.084922862e-13   pdiblc1 = -6.847759952e+00 lpdiblc1 = 2.173165875e-06 wpdiblc1 = 6.388363242e-06 ppdiblc1 = -1.913112088e-12   pdiblc2 = -1.639914392e-01 lpdiblc2 = 5.339842840e-08 wpdiblc2 = 1.496265006e-07 ppdiblc2 = -4.615705542e-14   pdiblcb = -5.425757567e+00 lpdiblcb = 1.763193186e-06 wpdiblcb = 4.328331535e-06 ppdiblcb = -1.474632506e-12   drout = 1.534104152e+01 ldrout = -4.539957100e-06 wdrout = -1.301520713e-05 pdrout = 3.978481657e-12   pscbe1 = 7.997817757e+08 lpscbe1 = 4.970591188e-02 wpscbe1 = 8.330606887e-02 ppscbe1 = -1.897492662e-8   pscbe2 = 5.377807903e-08 lpscbe2 = -1.236841807e-14 wpscbe2 = -3.197782513e-14 ppscbe2 = 8.716717985e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -1.934349062e+01 lbeta0 = 8.565588157e-06 wbeta0 = 2.394327047e-05 pbeta0 = -7.251069825e-12   agidl = 4.131073791e-09 lagidl = -9.002716537e-16 wagidl = -3.887613442e-15 pagidl = 8.946932164e-22   bgidl = 2.947568974e+09 lbgidl = -4.436076221e+02 wbgidl = -7.360195684e+02 pbgidl = 1.676469439e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.573018207e-01 lkt1 = -9.158349179e-08 wkt1 = -2.557326204e-07 pkt1 = 6.244087409e-14   kt2 = -1.817352677e+00 lkt2 = 5.248800270e-07 wkt2 = 1.517545794e-06 pkt2 = -4.514447169e-13   at = -4.985586615e+03 lat = 3.529920594e-02 wat = 1.270158479e-01 pat = -4.865039302e-8   ute = 2.282501354e+00 lute = -1.024506730e-06 wute = -4.514702832e-06 pute = 1.421054959e-12   ua1 = 1.818559352e-08 lua1 = -5.342422940e-15 wua1 = -1.540715798e-14 pua1 = 4.599859501e-21   ub1 = -2.937212874e-17 lub1 = 8.680664617e-24 wub1 = 2.403796889e-23 pub1 = -7.145802404e-30   uc1 = -1.426626737e-10 luc1 = -5.468405939e-18 wuc1 = -1.611171500e-16 puc1 = 6.294723428e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.98 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.6e-07 wmax = 9.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {3.995817037e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.025138049e-07 wvth0 = -1.224099744e-06 pvth0 = 2.527745365e-13   k1 = -1.241388840e+01 lk1 = 2.863732605e-06 wk1 = 1.079589779e-05 pk1 = -2.286847476e-12   k2 = 5.882635846e+00 lk2 = -1.291586644e-06 wk2 = -4.798997049e-06 pk2 = 1.011676852e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 6.229557890e+01 ldsub = -1.332202861e-05 wdsub = -4.934912245e-05 pdsub = 1.060596259e-11   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {2.805093316e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.725867328e-07 wvoff = -2.400742544e-06 pvoff = 5.320755647e-13   nfactor = {-2.131213862e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.474930296e-06 wnfactor = 1.896316971e-05 pnfactor = -3.651627103e-12   eta0 = 1.777960789e+01 leta0 = -3.793626928e-06 weta0 = -1.396731495e-05 peta0 = 3.017028571e-12   etab = 1.757363737e+00 letab = -3.634997767e-07 wetab = -1.434191271e-06 petab = 2.926441386e-13   u0 = -2.183709527e-01 lu0 = 4.538348704e-08 wu0 = 1.840740511e-07 pu0 = -3.752189218e-14   ua = -8.999059598e-08 lua = 1.772852943e-14 wua = 7.186493182e-14 pua = -1.434510943e-20   ub = 7.770823732e-17 lub = -1.518564252e-23 wub = -6.227383524e-23 pub = 1.231426540e-29   uc = -8.831804458e-10 luc = 1.896163089e-16 wuc = 7.033426684e-16 puc = -1.509927184e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.155471555e+06 lvsat = -9.442932567e-02 wvsat = -3.641680554e+00 pvsat = 7.565117766e-7   a0 = -9.253595110e+00 la0 = 1.958772635e-06 wa0 = 8.451759989e-06 pa0 = -1.604035167e-12   ags = 1.249999302e+00 lags = 1.500191296e-13 wags = 6.097528313e-13 pags = -1.309596627e-19   a1 = 0.0   a2 = -1.286221372e+01 la2 = 3.103383557e-06 wa2 = 1.062097850e-05 pa2 = -2.438198331e-12   b0 = 0.0   b1 = 0.0   keta = -4.562756898e+00 lketa = 9.785028387e-07 wketa = 3.634715933e-06 pketa = -7.793812187e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.116874927e+00 lpclm = -1.179956797e-06 wpclm = -4.375258987e-06 ppclm = 9.395499436e-13   pdiblc1 = 2.138352903e+01 lpdiblc1 = -4.574953527e-06 wpdiblc1 = -1.688055221e-05 ppdiblc1 = 3.639751464e-12   pdiblc2 = 5.899742714e-01 lpdiblc2 = -1.271681337e-07 wpdiblc2 = -4.658321081e-07 ppdiblc2 = 1.010468911e-13   pdiblcb = 1.984431253e+01 lpdiblcb = -4.290692200e-06 wpdiblcb = -1.613805969e-05 ppdiblcb = 3.424969126e-12   drout = -4.461562059e+01 ldrout = 9.797094913e-06 wdrout = 3.632061786e-05 pdrout = -7.800760702e-12   pscbe1 = 7.999999957e+08 lpscbe1 = 9.073963165e-07 wpscbe1 = 4.055702209e-06 ppscbe1 = -8.710632324e-13   pscbe2 = -9.720608779e-08 lpscbe2 = 2.366561378e-14 wpscbe2 = 8.247591043e-14 ppscbe2 = -1.864812240e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.431403522e+01 lbeta0 = -1.861563957e-05 wbeta0 = -6.834476244e-05 pbeta0 = 1.479754942e-11   agidl = 1.432703312e-09 lagidl = -3.069698457e-16 wagidl = 3.468248436e-16 pagidl = -7.501593629e-23   bgidl = 9.999964570e+08 lbgidl = 7.609389763e-04 wbgidl = 3.104705856e-03 pbgidl = -6.668132000e-10   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 5.344273521e-01 lkt1 = -2.677368392e-07 wkt1 = -8.275898344e-07 pkt1 = 2.070775018e-13   kt2 = 4.662866758e+00 lkt2 = -1.022141235e-06 wkt2 = -3.789368238e-06 pkt2 = 8.138615633e-13   at = 1.722814941e+06 lat = -3.849886100e-01 wat = -1.323117314e+00 pat = 3.026749269e-7   ute = -1.959926881e+01 lute = 4.255139445e-06 wute = 1.552835261e-05 pute = -3.378923420e-12   ua1 = -4.831595733e-08 lua1 = 1.053676213e-14 wua1 = 3.906277271e-14 pua1 = -8.389707011e-21   ub1 = 7.468287873e-17 lub1 = -1.614151794e-23 wub1 = -5.984119789e-23 pub1 = 1.285239328e-29   uc1 = -1.202828265e-09 luc1 = 2.536254920e-16 wuc1 = 9.402618090e-16 puc1 = -2.019447300e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.99 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.100 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.143767018e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.319531148e-07 wvth0 = 7.105427358e-21   k1 = 4.210177391e-01 lk1 = 2.132656424e-7   k2 = 5.626381206e-02 lk2 = -3.000267020e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 1.016439537e-26 pcit = 8.131516294e-32   voff = {-1.699412101e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.680610028e-7   nfactor = {1.682760886e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.726492433e-7   eta0 = 0.08   etab = -0.07   u0 = 6.320637964e-03 lu0 = 3.088464059e-8   ua = -7.269192156e-10 lua = 1.507603820e-16   ub = 1.320154755e-19 lub = 9.547120828e-24   uc = -1.283886196e-10 luc = 4.555983095e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.640088689e+04 lvsat = 1.077670413e+0   a0 = 1.632011387e+00 la0 = -3.368254479e-6   ags = 2.730837312e-04 lags = 2.265737709e-6   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 4.581250717e-08 lb0 = -3.686887499e-13   b1 = -6.681756343e-09 lb1 = 5.377327165e-14   keta = 4.028268441e-02 lketa = -3.392369294e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 wpclm = 1.110223025e-22 ppclm = -1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 1.919546137e-03 lpdiblc2 = -1.287843679e-8   pdiblcb = -2.718651916e-01 lpdiblcb = 9.395428170e-7   drout = 0.56   pscbe1 = 8.000326941e+08 lpscbe1 = -6.554436787e-1   pscbe2 = 1.316918687e-08 lpscbe2 = -6.231974900e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.590871467e+01 lbeta0 = -3.189343322e-4   agidl = 2.876157201e-09 lagidl = -1.956461964e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = -4.267601714e-01 legidl = 1.056036940e-05 wegidl = 8.881784197e-22 pegidl = 7.105427358e-27   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.365589613e-01 lkt1 = -3.390156381e-8   kt2 = -6.269565276e-02 lkt2 = 8.319130491e-8   at = 1.185992956e+05 lat = -9.544604462e-1   ute = -4.992636630e-02 lute = -6.626518113e-7   ua1 = 2.269582021e-09 lua1 = -3.596210395e-15   ub1 = -1.572949839e-18 lub1 = 6.897433758e-24   uc1 = -4.389120218e-11 luc1 = 2.827177762e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.101 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539359e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584525e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-08 ppdiblc2 = -1.387778781e-29   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+03 wpscbe1 = -7.629394531e-12   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901147e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-7   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23 pub1 = 2.465190329e-44   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.102 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308607e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = -5.551115123e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = 1.332267630e-21 ppclm = 6.217248938e-27   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16 wagidl = -1.654361225e-30   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343240e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-07 wute = -8.881784197e-22   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 wuc1 = 5.169878828e-32 puc1 = 1.033975766e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.103 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-08 wk2 = -2.220446049e-22 pk2 = 2.220446049e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-06 pdsub = 3.552713679e-27   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = 3.400058013e-22 peta0 = -2.428612866e-28   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = -4.787836794e-22 petab = -2.872702076e-27   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493533e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554777e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463397e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = 1.776356839e-21 pute = -5.329070518e-27   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24 wub1 = 1.232595164e-38   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 wuc1 = 4.135903063e-31 puc1 = -4.135903063e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.104 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140123256e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.326188593e-8   k1 = 5.232439484e-01 lk1 = -7.393371107e-9   k2 = -1.226088730e-02 lk2 = 2.100073728e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.277500803e+00 ldsub = -5.246443427e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.926698888e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.316212391e-9   nfactor = {1.185783805e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.894038578e-7   eta0 = -3.486985538e-02 leta0 = 2.670462627e-07 peta0 = 8.881784197e-28   etab = -1.729964684e+00 letab = 9.472731180e-7   u0 = 1.389723133e-02 lu0 = -4.306283297e-9   ua = -9.132162872e-10 lua = -1.574263421e-16   ub = 2.527606944e-18 lub = -7.074172299e-25   uc = -1.014940739e-10 luc = 3.852094380e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.311994564e+04 lvsat = 1.157790805e-1   a0 = 8.881460474e-01 la0 = -7.713305401e-8   ags = 1.120744391e-01 lags = 6.233271741e-7   a1 = 0.0   a2 = 1.053132798e+00 la2 = -5.568169504e-8   b0 = -9.608784530e-17 lb0 = 1.006784421e-22   b1 = -3.994811609e-20 lb1 = 4.185663734e-26   keta = 1.311717861e-02 lketa = -2.809313044e-08 pketa = -5.551115123e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.624337286e+00 lpclm = -8.573312648e-7   pdiblc1 = 6.467424655e-02 lpdiblc1 = -2.690083368e-8   pdiblc2 = 7.922616047e-04 lpdiblc2 = -3.795686529e-10   pdiblcb = -1.354002314e-02 lpdiblcb = -1.200747726e-8   drout = 1.041454917e+00 ldrout = -4.343542515e-8   pscbe1 = 8.275046100e+08 lpscbe1 = -4.317079225e+1   pscbe2 = 3.162763138e-09 lpscbe2 = 6.301310952e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.507657499e+00 lbeta0 = 1.216018119e-6   agidl = 1.064658721e-09 lagidl = -5.831934307e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.190246567e-01 lkt1 = -6.290849829e-8   kt2 = -6.368883441e-02 lkt2 = 1.585247260e-8   at = 8.716611382e+04 lat = -2.661806463e-02 wat = 4.656612873e-16   ute = -1.975547800e+00 lute = 9.716939615e-7   ua1 = -3.637135874e-09 lua1 = 3.359933500e-15 wua1 = 3.308722450e-30 pua1 = -3.308722450e-36   ub1 = 4.413339682e-18 lub1 = -3.686548278e-24 pub1 = 6.162975822e-45   uc1 = 3.433541843e-10 luc1 = -2.896421036e-16 puc1 = 4.135903063e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.105 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.083758130e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.386478892e-9   k1 = 4.286126363e-01 lk1 = 4.444329585e-8   k2 = 2.077621672e-02 lk2 = -1.599682593e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.339715233e-01 ldsub = 3.033024110e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.158159998e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.362648555e-9   nfactor = {1.886976015e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.053082948e-7   eta0 = 4.081427101e-01 leta0 = 2.437505465e-8   etab = -1.347621329e-03 letab = 3.799063485e-10   u0 = 7.040683625e-03 lu0 = -5.504378792e-10   ua = -1.613983779e-09 lua = 2.264365708e-16   ub = 2.025147933e-18 lub = -4.321827452e-25   uc = -6.712093967e-11 luc = 1.969220019e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.716932025e+05 lvsat = -1.284569167e-2   a0 = 9.052648244e-01 la0 = -8.651029208e-8   ags = 9.445453886e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.136650759e+00 la2 = -1.014307462e-7   b0 = 1.921756906e-16 lb0 = -5.722511627e-23   b1 = 7.989623218e-20 lb1 = -2.379110054e-26   keta = -4.583734636e-02 lketa = 4.200684472e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.292099820e-01 lpclm = 3.771055897e-07 ppclm = -2.220446049e-28   pdiblc1 = -4.478501477e-01 lpdiblc1 = 2.538472164e-07 wpdiblc1 = -4.440892099e-22 ppdiblc1 = 3.330669074e-28   pdiblc2 = -9.997833428e-03 lpdiblc2 = 5.530975654e-09 wpdiblc2 = 3.469446952e-24 ppdiblc2 = -9.974659987e-30   pdiblcb = 2.653629919e-01 lpdiblcb = -1.647835763e-07 wpdiblcb = -4.440892099e-22 ppdiblcb = -2.220446049e-28   drout = 1.478478000e+00 ldrout = -2.828257447e-7   pscbe1 = 6.876139896e+08 lpscbe1 = 3.345779234e+1   pscbe2 = 2.160022972e-08 lpscbe2 = -3.798272305e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.510363785e+00 lbeta0 = 1.189856830e-7   agidl = 1.490566362e-12 lagidl = -8.164949889e-19   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.471888216e-01 lkt1 = 7.296627166e-9   kt2 = -1.323292858e-02 lkt2 = -1.178601122e-8   at = 3.656378506e+03 lat = 1.912648063e-2   ute = 5.522314189e-01 lute = -4.129603001e-7   ua1 = 5.118987964e-09 lua1 = -1.436452236e-15 pua1 = 6.617444900e-36   ub1 = -4.874445755e-18 lub1 = 1.401068390e-24   uc1 = -2.896530271e-10 luc1 = 5.710342159e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.106 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.072602848e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.352851598e-10   k1 = -1.155995736e+00 lk1 = 5.163000540e-7   k2 = 6.092877219e-01 lk2 = -1.912408394e-07 pk2 = -4.440892099e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.329682527e+00 ldsub = -4.600896739e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.145411686e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.579446431e-8   nfactor = {2.861935894e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.850103831e-7   eta0 = 1.370249058e+00 leta0 = -2.621161630e-07 peta0 = -1.776356839e-27   etab = 8.874965423e-02 letab = -2.644880988e-08 wetab = -1.457167720e-22 petab = -2.645453301e-29   u0 = 3.544653257e-03 lu0 = 4.905925638e-10   ua = -6.707151893e-10 lua = -5.444523355e-17   ub = 3.530366730e-19 lub = 6.573018533e-26   uc = -4.489843184e-12 luc = 1.042225433e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.942483259e+05 lvsat = -4.933954354e-2   a0 = -1.072606605e+00 la0 = 5.024503727e-7   ags = 2.340909298e+00 lags = -2.484818634e-7   a1 = 0.0   a2 = 1.286764451e+00 la2 = -1.461308507e-7   b0 = 0.0   b1 = 0.0   keta = -1.374979945e-01 lketa = 3.149493397e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.864146677e-01 lpclm = -1.465454032e-8   pdiblc1 = 1.175483577e+00 lpdiblc1 = -2.295409836e-7   pdiblc2 = 2.392678142e-02 lpdiblc2 = -4.570926532e-9   pdiblcb = 1.026049661e-02 lpdiblcb = -8.882043078e-8   drout = -1.004957054e+00 ldrout = 4.566791284e-7   pscbe1 = 7.998864011e+08 lpscbe1 = 2.587501007e-2   pscbe2 = 1.361663723e-08 lpscbe2 = -1.420958051e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.072723056e+01 lbeta0 = -5.411418223e-7   agidl = -7.514396508e-10 lagidl = 2.233873004e-16 wagidl = -1.525114254e-30 pagidl = -4.135903063e-37   bgidl = 2.023190692e+09 lbgidl = -2.330572500e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.784803471e-01 lkt1 = -1.316303884e-8   kt2 = 8.855639745e-02 lkt2 = -4.209632778e-8   at = 1.545355679e+05 lat = -2.580156999e-2   ute = -3.387583285e+00 lute = 7.602180233e-7   ua1 = -1.164492862e-09 lua1 = 4.346112672e-16   ub1 = 8.175256375e-19 lub1 = -2.938583918e-25 pub1 = 7.703719778e-46   uc1 = -3.450121774e-10 luc1 = 7.358799255e-17 wuc1 = 1.654361225e-30   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.107 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 8.6e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-3.508192265e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.951663093e-07 wvth0 = 1.887394939e-06 pvth0 = -4.619870962e-13   k1 = 2.469509058e+00 lk1 = -3.325987984e-07 wk1 = -1.054739539e-06 pk1 = 2.581738707e-13   k2 = 3.186247087e+00 lk2 = -8.362893388e-07 wk2 = -2.652046034e-06 pk2 = 6.491545681e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 6.086699853e-01 ldsub = -7.316764778e-08 wdsub = -2.320315973e-07 pdsub = 5.679553423e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {4.788801034e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.729743274e-07 wvoff = -5.485371461e-07 pvoff = 1.342681799e-13   nfactor = {2.013653175e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.427207843e-06 wnfactor = -1.403958799e-05 pnfactor = 3.436540151e-12   eta0 = 9.504626002e-01 leta0 = -1.789259875e-07 weta0 = -5.674109380e-07 peta0 = 1.388880124e-13   etab = -6.838737668e-01 letab = 1.606960796e-07 wetab = 5.096001490e-07 petab = -1.247373765e-13   u0 = 2.888374633e-01 lu0 = -6.930533960e-08 wu0 = -2.197815203e-07 pu0 = 5.379702164e-14   ua = 4.588435905e-08 lua = -1.145402705e-14 wua = -3.632305537e-14 pua = 8.890975879e-21   ub = -4.490443391e-17 lub = 1.114853332e-23 wub = 3.535429720e-23 pub = -8.653848097e-30   uc = 2.975000542e-12 luc = -7.071951356e-19 wuc = -2.242654996e-18 puc = 5.489458766e-25   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.390959344e+08 lvsat = 3.406620996e+01 wvsat = 1.080309769e+02 pvsat = -2.644328237e-5   a0 = 1.020239189e+01 la0 = -2.219886972e-06 wa0 = -7.039719452e-06 pa0 = 1.723147329e-12   ags = 1.249999979e+00 lags = 7.332786822e-15 wags = 7.087425047e-14 pags = -1.734824195e-20   a1 = 0.0   a2 = -6.057881237e+00 la2 = 1.640748313e-06 wa2 = 5.203151242e-06 pa2 = -1.273601345e-12   b0 = 0.0   b1 = 0.0   keta = 5.509224699e-02 lketa = -1.329571621e-08 wketa = -4.216332680e-08 pketa = 1.032052832e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.158332438e-01 lpclm = 1.528285266e-09 wpclm = 4.846434589e-09 ppclm = -1.186286027e-15   pdiblc1 = 7.750135355e-01 lpdiblc1 = -1.486477334e-07 wpdiblc1 = -4.713927041e-07 ppdiblc1 = 1.153851492e-13   pdiblc2 = 4.643887972e-02 lpdiblc2 = -1.042247675e-08 wpdiblc2 = -3.305183604e-08 ppdiblc2 = 8.090263166e-15   pdiblcb = -2.132836524e+00 lpdiblcb = 4.291270246e-07 wpdiblcb = 1.360849654e-06 ppdiblcb = -3.331019742e-13   drout = 1.000002816e+00 ldrout = -6.510571069e-13 wdrout = -1.198092463e-12 pdrout = 2.932630778e-19   pscbe1 = 8.000000146e+08 lpscbe1 = -3.551727295e-06 wpscbe1 = -1.094653320e-05 ppscbe1 = 2.679435730e-12   pscbe2 = -3.249434666e-08 lpscbe2 = 9.759804745e-15 wpscbe2 = 3.095035136e-14 ppscbe2 = -7.575872255e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.342122330e+01 lbeta0 = -1.240952045e-06 wbeta0 = -3.935317022e-06 pbeta0 = 9.632672240e-13   agidl = 6.548006742e-08 lagidl = -1.597175732e-14 wagidl = -5.064973598e-14 pagidl = 1.239778912e-20   bgidl = 1.000000366e+09 lbgidl = -7.891886902e-05 wbgidl = -7.796936035e-06 pbgidl = 1.908493042e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 7.104138873e-01 lkt1 = -3.051570492e-07 wkt1 = -9.677159453e-07 pkt1 = 2.368726705e-13   kt2 = -9.625899383e-02 lkt2 = -2.176820502e-15 wkt2 = -2.204999205e-14 pkt2 = 5.397287950e-21   at = 8.308254398e+05 lat = -1.932661250e-01 wat = -6.128867295e-01 pat = 1.500193492e-7   ute = -1.920026367e+00 lute = 4.577356939e-07 wute = 1.451574046e-06 pute = -3.553090372e-13   ua1 = 7.435795451e-10 lua1 = 8.034989610e-23 wua1 = -4.491645519e-22 pua1 = 1.099442545e-28   ub1 = -4.726033506e-19 lub1 = 7.935641432e-31 wub1 = 1.912867566e-30 pub1 = -4.682221595e-37   uc1 = -2.193904617e-11 luc1 = 1.085018434e-23 wuc1 = 2.417686390e-23 puc1 = -5.917891639e-30   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.108 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.109 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.143767018e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.319531148e-7   k1 = 4.210177391e-01 lk1 = 2.132656424e-7   k2 = 5.626381206e-02 lk2 = -3.000267020e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 6.776263578e-27 pcit = -1.355252716e-31   voff = {-1.699412101e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.680610028e-7   nfactor = {1.682760886e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.726492433e-7   eta0 = 0.08   etab = -0.07   u0 = 6.320637964e-03 lu0 = 3.088464059e-8   ua = -7.269192156e-10 lua = 1.507603820e-16   ub = 1.320154755e-19 lub = 9.547120828e-24   uc = -1.283886196e-10 luc = 4.555983095e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.640088689e+04 lvsat = 1.077670413e+0   a0 = 1.632011387e+00 la0 = -3.368254479e-6   ags = 2.730837313e-04 lags = 2.265737709e-6   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 4.581250717e-08 lb0 = -3.686887499e-13   b1 = -6.681756343e-09 lb1 = 5.377327165e-14   keta = 4.028268441e-02 lketa = -3.392369294e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 ppclm = 1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 1.919546137e-03 lpdiblc2 = -1.287843679e-8   pdiblcb = -2.718651916e-01 lpdiblcb = 9.395428170e-7   drout = 0.56   pscbe1 = 8.000326941e+08 lpscbe1 = -6.554436786e-1   pscbe2 = 1.316918687e-08 lpscbe2 = -6.231974900e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.590871467e+01 lbeta0 = -3.189343322e-4   agidl = 2.876157201e-09 lagidl = -1.956461964e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = -4.267601714e-01 legidl = 1.056036940e-05 pegidl = -2.842170943e-26   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.365589613e-01 lkt1 = -3.390156381e-8   kt2 = -6.269565276e-02 lkt2 = 8.319130491e-8   at = 1.185992956e+05 lat = -9.544604462e-1   ute = -4.992636630e-02 lute = -6.626518113e-7   ua1 = 2.269582021e-09 lua1 = -3.596210395e-15   ub1 = -1.572949839e-18 lub1 = 6.897433758e-24   uc1 = -4.389120218e-11 luc1 = 2.827177762e-16 puc1 = -1.654361225e-36   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.110 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539359e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584524e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-08 ppdiblc2 = -1.387778781e-29   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 ppscbe2 = 4.235164736e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-7   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.111 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308607e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = -8.881784197e-22 ppclm = 2.664535259e-27   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343240e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.112 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-08 wk2 = 2.220446049e-22 pk2 = 2.220446049e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-06 pdsub = 3.552713679e-27   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-07 wnfactor = 1.421085472e-20   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = 3.573530361e-22 peta0 = -8.326672685e-29   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = -4.510281038e-22 petab = 3.053113318e-28   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493533e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554778e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463397e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = -8.881784197e-22   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24 wub1 = 1.232595164e-38 pub1 = 1.232595164e-44   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 wuc1 = -2.067951531e-31 puc1 = -4.135903063e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.113 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140123256e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.326188593e-8   k1 = 5.232439484e-01 lk1 = -7.393371107e-9   k2 = -1.226088730e-02 lk2 = 2.100073728e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.277500803e+00 ldsub = -5.246443427e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.926698888e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.316212391e-9   nfactor = {1.185783805e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.894038578e-7   eta0 = -3.486985538e-02 leta0 = 2.670462627e-7   etab = -1.729964684e+00 letab = 9.472731180e-7   u0 = 1.389723133e-02 lu0 = -4.306283297e-9   ua = -9.132162872e-10 lua = -1.574263421e-16   ub = 2.527606944e-18 lub = -7.074172299e-25   uc = -1.014940739e-10 luc = 3.852094380e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.311994564e+04 lvsat = 1.157790805e-01 pvsat = 2.328306437e-22   a0 = 8.881460474e-01 la0 = -7.713305401e-8   ags = 1.120744391e-01 lags = 6.233271741e-7   a1 = 0.0   a2 = 1.053132798e+00 la2 = -5.568169504e-8   b0 = -9.608784530e-17 lb0 = 1.006784421e-22   b1 = -3.994811609e-20 lb1 = 4.185663734e-26   keta = 1.311717861e-02 lketa = -2.809313044e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.624337286e+00 lpclm = -8.573312648e-7   pdiblc1 = 6.467424655e-02 lpdiblc1 = -2.690083368e-8   pdiblc2 = 7.922616047e-04 lpdiblc2 = -3.795686529e-10   pdiblcb = -1.354002314e-02 lpdiblcb = -1.200747726e-8   drout = 1.041454917e+00 ldrout = -4.343542515e-8   pscbe1 = 8.275046100e+08 lpscbe1 = -4.317079225e+1   pscbe2 = 3.162763138e-09 lpscbe2 = 6.301310952e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.507657499e+00 lbeta0 = 1.216018119e-6   agidl = 1.064658721e-09 lagidl = -5.831934307e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.190246567e-01 lkt1 = -6.290849829e-8   kt2 = -6.368883441e-02 lkt2 = 1.585247260e-8   at = 8.716611382e+04 lat = -2.661806463e-2   ute = -1.975547800e+00 lute = 9.716939615e-7   ua1 = -3.637135874e-09 lua1 = 3.359933500e-15 wua1 = 6.617444900e-30 pua1 = 1.654361225e-36   ub1 = 4.413339682e-18 lub1 = -3.686548278e-24 wub1 = -1.232595164e-38   uc1 = 3.433541843e-10 luc1 = -2.896421036e-16 wuc1 = -8.271806126e-31 puc1 = 8.271806126e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.114 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.083758130e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.386478892e-9   k1 = 4.286126363e-01 lk1 = 4.444329585e-8   k2 = 2.077621672e-02 lk2 = -1.599682593e-08 pk2 = -2.775557562e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.339715233e-01 ldsub = 3.033024110e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.158159998e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.362648555e-9   nfactor = {1.886976015e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.053082948e-7   eta0 = 4.081427101e-01 leta0 = 2.437505465e-8   etab = -1.347621329e-03 letab = 3.799063485e-10   u0 = 7.040683625e-03 lu0 = -5.504378792e-10   ua = -1.613983779e-09 lua = 2.264365708e-16   ub = 2.025147933e-18 lub = -4.321827452e-25 wub = 1.232595164e-38   uc = -6.712093967e-11 luc = 1.969220019e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.716932025e+05 lvsat = -1.284569167e-2   a0 = 9.052648244e-01 la0 = -8.651029208e-8   ags = 9.445453886e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.136650759e+00 la2 = -1.014307462e-7   b0 = 1.921756906e-16 lb0 = -5.722511627e-23   b1 = 7.989623218e-20 lb1 = -2.379110054e-26   keta = -4.583734636e-02 lketa = 4.200684472e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.292099820e-01 lpclm = 3.771055897e-07 wpclm = 8.881784197e-22 ppclm = -6.661338148e-28   pdiblc1 = -4.478501477e-01 lpdiblc1 = 2.538472164e-07 wpdiblc1 = 4.440892099e-22 ppdiblc1 = -2.775557562e-28   pdiblc2 = -9.997833428e-03 lpdiblc2 = 5.530975654e-09 wpdiblc2 = 1.821459650e-23 ppdiblc2 = 5.854691731e-30   pdiblcb = 2.653629919e-01 lpdiblcb = -1.647835763e-07 wpdiblcb = -4.440892099e-22 ppdiblcb = -1.110223025e-28   drout = 1.478478000e+00 ldrout = -2.828257447e-7   pscbe1 = 6.876139896e+08 lpscbe1 = 3.345779234e+1   pscbe2 = 2.160022972e-08 lpscbe2 = -3.798272305e-15 wpscbe2 = -1.058791184e-28   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.510363785e+00 lbeta0 = 1.189856830e-7   agidl = 1.490566362e-12 lagidl = -8.164949889e-19   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.471888216e-01 lkt1 = 7.296627166e-9   kt2 = -1.323292858e-02 lkt2 = -1.178601122e-8   at = 3.656378506e+03 lat = 1.912648063e-2   ute = 5.522314189e-01 lute = -4.129603001e-07 pute = -4.440892099e-28   ua1 = 5.118987964e-09 lua1 = -1.436452236e-15   ub1 = -4.874445755e-18 lub1 = 1.401068390e-24   uc1 = -2.896530271e-10 luc1 = 5.710342159e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.115 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-2.687610411e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.402992793e-07 wvth0 = -6.239677336e-07 pvth0 = 1.858019919e-13   k1 = -1.528203460e+00 lk1 = 6.271342089e-07 wk1 = 2.889195456e-07 pk1 = -8.603301769e-14   k2 = 9.039665489e-02 lk2 = -3.672805190e-08 wk2 = 4.027798507e-07 pk2 = -1.199377701e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 3.514802141e+00 ldsub = -8.129886668e-07 wdsub = -9.199277678e-07 pdsub = 2.739314911e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {3.103268022e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.914271713e-08 wvoff = -1.129990798e-07 pvoff = 3.364830099e-14   nfactor = {-2.544375839e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.424854093e-06 wnfactor = 4.196552169e-06 pnfactor = -1.249628322e-12   eta0 = 3.906387132e+00 leta0 = -1.017314678e-06 weta0 = -1.968631530e-06 peta0 = 5.862092538e-13   etab = 3.417117197e-01 letab = -1.017745889e-07 wetab = -1.963572500e-07 petab = 5.847028012e-14   u0 = -9.319903870e-02 lu0 = 2.929844544e-08 wu0 = 7.509554950e-08 pu0 = -2.236157725e-14   ua = -1.274241846e-08 lua = 3.540206207e-15 wua = 9.370442370e-15 pua = -2.790283477e-21   ub = 1.065501668e-17 lub = -3.001941910e-24 wub = -7.996726543e-24 pub = 2.381225246e-30   uc = -1.324958591e-10 luc = 3.915921681e-17 wuc = 9.936236572e-17 puc = -2.958762845e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.312455687e+07 lvsat = -3.869884671e+00 wvsat = -9.959296064e+00 pvsat = 2.965629385e-6   a0 = -3.474221113e+00 la0 = 1.217591133e-06 wa0 = 1.864210033e-06 pa0 = -5.551151425e-13   ags = 2.340909330e+00 lags = -2.484818730e-07 wags = -2.498975959e-14 pags = 7.441322225e-21   a1 = 0.0   a2 = 2.274002596e+00 la2 = -4.401056894e-07 wa2 = -7.663258401e-07 pa2 = 2.281926770e-13   b0 = 0.0   b1 = 0.0   keta = -2.624691141e-01 lketa = 6.870820910e-08 wketa = 9.700658208e-08 pketa = -2.888613498e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.739663685e-01 lpclm = -1.094774802e-08 wpclm = 9.662768204e-09 ppclm = -2.877330802e-15   pdiblc1 = 2.962673019e+00 lpdiblc1 = -7.617213196e-07 wpdiblc1 = -1.387273635e-06 ppdiblc1 = 4.130954065e-13   pdiblc2 = -1.085659118e-03 lpdiblc2 = 2.877152948e-09 wpdiblc2 = 1.941545674e-08 ppdiblc2 = -5.781437631e-15   pdiblcb = -7.233950901e+00 lpdiblcb = 2.068324618e-06 wpdiblcb = 5.623188702e-06 ppdiblcb = -1.674445016e-12   drout = -1.004958507e+00 ldrout = 4.566795611e-07 wdrout = 1.127828043e-12 pdrout = -3.358389939e-19   pscbe1 = 7.998864054e+08 lpscbe1 = 2.587371421e-02 wpscbe1 = -3.378005981e-06 ppscbe1 = 1.005886078e-12   pscbe2 = -7.596283286e-09 lpscbe2 = 4.895719355e-15 wpscbe2 = 1.646614772e-14 ppscbe2 = -4.903207137e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.075097328e+01 lbeta0 = -5.482118102e-07 wbeta0 = -1.842985752e-08 pbeta0 = 5.487950823e-15   agidl = -2.909597292e-08 lagidl = 8.663680694e-15 wagidl = 2.200193375e-14 pagidl = -6.551625821e-21   bgidl = 2.023190708e+09 lbgidl = -2.330572548e+02 wbgidl = -1.253784180e-05 pbgidl = 3.733459473e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -9.511726902e-01 lkt1 = 1.275929236e-07 wkt1 = 3.669189229e-07 pkt1 = -1.092592823e-13   kt2 = 5.223550138e-01 lkt2 = -1.712707108e-07 wkt2 = -3.367283676e-07 pkt2 = 1.002692897e-13   at = -6.467721351e+04 lat = 3.947451599e-02 wat = 1.701599757e-01 pat = -5.066938677e-8   ute = -7.520659927e+00 lute = 1.990944920e-06 wute = 3.208226348e-06 pute = -9.553296008e-13   ua1 = -4.919317356e-09 lua1 = 1.552704131e-15 wua1 = 2.914614927e-15 pua1 = -8.678994598e-22   ub1 = 4.239703480e-18 lub1 = -1.312897399e-24 wub1 = -2.656403951e-24 pub1 = 7.910106865e-31   uc1 = -4.152434317e-10 luc1 = 9.450110432e-17 wuc1 = 5.451574704e-17 puc1 = -1.623342657e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.116 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.2e-07 wmax = 8.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.617044431e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.179203723e-08 wvth0 = 4.194254735e-07 pvth0 = -5.572723822e-14   k1 = 1.225104074e+00 lk1 = -4.455661866e-13 wk1 = -8.879256905e-08 pk1 = 3.860341735e-19   k2 = -2.455172839e+00 lk2 = 5.836225208e-07 wk2 = 1.727004638e-06 pk2 = -4.530264546e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.446830879e-02 ldsub = 2.052340093e-12 wdsub = 2.827175669e-07 pdsub = -1.128433690e-18   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.725243638e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.229685509e-14 wvoff = 3.472704625e-08 pvoff = -1.866861687e-20   nfactor = {3.711166594e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.240142692e-12 wnfactor = -1.289693951e-06 pnfactor = 1.491454938e-18   eta0 = -5.599256183e-01 leta0 = -3.131386705e-13 weta0 = 6.050007296e-07 peta0 = 1.783030452e-19   etab = -1.051100985e-01 letab = 2.694352315e-13 wetab = 6.034526925e-08 petab = -1.463671004e-19   u0 = 8.197491316e-03 lu0 = 6.665800933e-09 wu0 = -1.939793637e-09 pu0 = -5.174208718e-15   ua = 2.801447964e-09 lua = -3.202058920e-19 wua = -2.880721134e-15 pua = 2.421050294e-25   ub = -2.524405275e-18 lub = 9.937095441e-31 wub = 2.457562815e-24 pub = -5.503894369e-37   uc = 3.942475727e-11 luc = -1.690401188e-24 wuc = -3.053612256e-17 puc = -3.057387410e-31   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.882216608e+07 lvsat = -2.268759603e+01 wvsat = -6.888634606e+01 pvsat = 1.761083796e-5   a0 = 1.871361671e+00 la0 = 1.089890716e-12 wa0 = -5.729072035e-07 pa0 = -8.210495039e-19   ags = 1.249999992e+00 lags = 1.604945510e-15 wags = 6.038987976e-14 pags = -1.290210605e-20   a1 = 0.0   a2 = 3.418077866e-01 la2 = -1.799187999e-14 wa2 = 2.355078315e-07 pa2 = 1.340958988e-20   b0 = 0.0   b1 = 0.0   keta = 3.918087929e-02 lketa = -1.269545023e-13 wketa = -2.981241403e-08 pketa = 6.647856664e-20   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.259020748e-01 lpclm = 1.036818915e-13 wpclm = -2.969314199e-09 ppclm = -6.257883811e-20   pdiblc1 = -3.815119025e-01 lpdiblc1 = 4.308279760e-13 wpdiblc1 = 4.263393497e-07 ppdiblc1 = -3.126736949e-19   pdiblc2 = 1.154586025e-02 lpdiblc2 = 9.267316692e-15 wpdiblc2 = -5.966757754e-09 ppdiblc2 = -4.002454618e-21   pdiblcb = 1.846606249e+00 lpdiblcb = 7.664284922e-13 wpdiblcb = -1.728121169e-06 ppdiblcb = -4.405485541e-19   drout = 1.000004799e+00 ldrout = -1.027174804e-12 wdrout = -2.737444305e-12 pdrout = 5.852176912e-19   pscbe1 = 7.999999844e+08 lpscbe1 = 3.500518799e-06 wpscbe1 = 1.245578003e-05 ppscbe1 = -2.794746399e-12   pscbe2 = 1.389738118e-08 lpscbe2 = -7.303075720e-23 wpscbe2 = -5.060392316e-15 ppscbe2 = 5.582279053e-28   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.344152637e+00 lbeta0 = 1.893961553e-12 wbeta0 = 5.667694638e-09 pbeta0 = -9.339867120e-19   agidl = 8.940163103e-09 lagidl = -2.021947716e-22 wagidl = -6.761652967e-15 pagidl = 1.529061560e-28   bgidl = 1.000000390e+09 lbgidl = -8.599177551e-05 wbgidl = -2.637344360e-05 pbgidl = 7.398712158e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.910009998e-01 lkt1 = -1.968219578e-13 wkt1 = -1.127624647e-07 pkt1 = 1.566699623e-19   kt2 = -2.295736492e-01 lkt2 = -1.714585425e-13 wkt2 = 1.034830795e-07 pkt2 = 1.367991773e-19   at = 1.086275108e+05 lat = 3.481948795e-08 wat = -5.229358668e-02 pat = -2.858058549e-14   ute = 1.220180155e+00 lute = 7.598353768e-14 wute = -9.859547429e-07 pute = -2.996962678e-21   ua1 = 1.897508409e-09 lua1 = 1.764838290e-21 wua1 = -8.957169594e-16 pua1 = -1.197609541e-27   ub1 = -1.524307226e-18 lub1 = 1.501840664e-31 wub1 = 8.163681156e-25 pub1 = 3.119004718e-38   uc1 = -3.555859511e-13 luc1 = 2.713569370e-23 wuc1 = -1.675374831e-17 puc1 = -1.855922558e-29   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.117 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.118 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.143767018e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.319531148e-7   k1 = 4.210177391e-01 lk1 = 2.132656424e-7   k2 = 5.626381206e-02 lk2 = -3.000267020e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 pcit = 1.490777987e-31   voff = {-1.699412101e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.680610028e-7   nfactor = {1.682760886e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.726492433e-7   eta0 = 0.08   etab = -0.07   u0 = 6.320637964e-03 lu0 = 3.088464059e-8   ua = -7.269192156e-10 lua = 1.507603820e-16   ub = 1.320154755e-19 lub = 9.547120828e-24   uc = -1.283886196e-10 luc = 4.555983095e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.640088689e+04 lvsat = 1.077670413e+0   a0 = 1.632011387e+00 la0 = -3.368254479e-6   ags = 2.730837313e-04 lags = 2.265737709e-06 pags = -3.552713679e-27   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-06 wa2 = -3.552713679e-21   b0 = 4.581250717e-08 lb0 = -3.686887499e-13   b1 = -6.681756343e-09 lb1 = 5.377327165e-14   keta = 4.028268441e-02 lketa = -3.392369294e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-6   pdiblc1 = 0.39   pdiblc2 = 1.919546137e-03 lpdiblc2 = -1.287843679e-8   pdiblcb = -2.718651916e-01 lpdiblcb = 9.395428170e-07 wpdiblcb = 8.881784197e-22   drout = 0.56   pscbe1 = 8.000326941e+08 lpscbe1 = -6.554436787e-1   pscbe2 = 1.316918687e-08 lpscbe2 = -6.231974900e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.590871467e+01 lbeta0 = -3.189343322e-04 pbeta0 = 9.094947018e-25   agidl = 2.876157201e-09 lagidl = -1.956461964e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = -4.267601714e-01 legidl = 1.056036940e-05 pegidl = -7.105427358e-27   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.365589613e-01 lkt1 = -3.390156381e-8   kt2 = -6.269565276e-02 lkt2 = 8.319130491e-8   at = 1.185992956e+05 lat = -9.544604462e-1   ute = -4.992636630e-02 lute = -6.626518113e-7   ua1 = 2.269582021e-09 lua1 = -3.596210395e-15   ub1 = -1.572949839e-18 lub1 = 6.897433758e-24   uc1 = -4.389120218e-11 luc1 = 2.827177762e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.119 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539358e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584525e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-08 wpdiblc2 = 1.734723476e-24   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 ppscbe2 = 1.058791184e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-7   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23 pub1 = -2.465190329e-44   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.120 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-08 wvoff = -8.881784197e-22   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308608e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = 5.551115123e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = -6.661338148e-22 ppclm = 1.332267630e-27   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343240e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 wuc1 = -2.584939414e-32 puc1 = -5.169878828e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.121 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-08 pk2 = -1.110223025e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = 1.353084311e-22 peta0 = -4.787836794e-28   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = 1.283695372e-22 petab = 2.706168623e-27   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-02 wvsat = -2.328306437e-16   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493534e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554778e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463397e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 pute = -3.552713679e-27   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 wuc1 = 2.067951531e-31 puc1 = -2.067951531e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.122 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140123256e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.326188593e-8   k1 = 5.232439484e-01 lk1 = -7.393371107e-9   k2 = -1.226088730e-02 lk2 = 2.100073728e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.277500803e+00 ldsub = -5.246443427e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.926698888e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.316212391e-9   nfactor = {1.185783805e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.894038578e-7   eta0 = -3.486985538e-02 leta0 = 2.670462627e-7   etab = -1.729964684e+00 letab = 9.472731180e-7   u0 = 1.389723133e-02 lu0 = -4.306283297e-9   ua = -9.132162872e-10 lua = -1.574263421e-16   ub = 2.527606944e-18 lub = -7.074172299e-25   uc = -1.014940739e-10 luc = 3.852094380e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.311994564e+04 lvsat = 1.157790805e-01 pvsat = -1.164153218e-22   a0 = 8.881460474e-01 la0 = -7.713305401e-08 wa0 = 3.552713679e-21   ags = 1.120744391e-01 lags = 6.233271741e-7   a1 = 0.0   a2 = 1.053132798e+00 la2 = -5.568169504e-8   b0 = -9.608784530e-17 lb0 = 1.006784421e-22   b1 = -3.994811609e-20 lb1 = 4.185663734e-26   keta = 1.311717861e-02 lketa = -2.809313044e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.624337286e+00 lpclm = -8.573312648e-7   pdiblc1 = 6.467424655e-02 lpdiblc1 = -2.690083368e-08 wpdiblc1 = -2.220446049e-22   pdiblc2 = 7.922616047e-04 lpdiblc2 = -3.795686529e-10   pdiblcb = -1.354002314e-02 lpdiblcb = -1.200747726e-8   drout = 1.041454917e+00 ldrout = -4.343542515e-8   pscbe1 = 8.275046100e+08 lpscbe1 = -4.317079225e+1   pscbe2 = 3.162763138e-09 lpscbe2 = 6.301310952e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.507657499e+00 lbeta0 = 1.216018119e-6   agidl = 1.064658721e-09 lagidl = -5.831934307e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.190246567e-01 lkt1 = -6.290849829e-8   kt2 = -6.368883441e-02 lkt2 = 1.585247260e-8   at = 8.716611382e+04 lat = -2.661806463e-2   ute = -1.975547800e+00 lute = 9.716939615e-7   ua1 = -3.637135874e-09 lua1 = 3.359933500e-15 wua1 = 3.308722450e-30 pua1 = 3.308722450e-36   ub1 = 4.413339682e-18 lub1 = -3.686548278e-24 pub1 = 6.162975822e-45   uc1 = 3.433541843e-10 luc1 = -2.896421036e-16 wuc1 = 4.135903063e-31   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.123 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.083758130e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.386478892e-9   k1 = 4.286126363e-01 lk1 = 4.444329585e-8   k2 = 2.077621672e-02 lk2 = -1.599682593e-08 pk2 = 2.775557562e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.339715233e-01 ldsub = 3.033024110e-07 pdsub = 4.440892099e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.158159998e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.362648555e-9   nfactor = {1.886976015e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.053082948e-7   eta0 = 4.081427101e-01 leta0 = 2.437505465e-8   etab = -1.347621329e-03 letab = 3.799063485e-10   u0 = 7.040683625e-03 lu0 = -5.504378792e-10   ua = -1.613983779e-09 lua = 2.264365708e-16   ub = 2.025147933e-18 lub = -4.321827452e-25   uc = -6.712093967e-11 luc = 1.969220019e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.716932025e+05 lvsat = -1.284569167e-2   a0 = 9.052648244e-01 la0 = -8.651029208e-8   ags = 9.445453886e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.136650759e+00 la2 = -1.014307462e-7   b0 = 1.921756906e-16 lb0 = -5.722511627e-23   b1 = 7.989623218e-20 lb1 = -2.379110054e-26   keta = -4.583734636e-02 lketa = 4.200684472e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.292099820e-01 lpclm = 3.771055897e-07 wpclm = 4.440892099e-22 ppclm = 1.110223025e-28   pdiblc1 = -4.478501477e-01 lpdiblc1 = 2.538472164e-07 wpdiblc1 = 7.771561172e-22 ppdiblc1 = 3.053113318e-28   pdiblc2 = -9.997833428e-03 lpdiblc2 = 5.530975654e-09 wpdiblc2 = 6.071532166e-24 ppdiblc2 = -1.084202172e-30   pdiblcb = 2.653629919e-01 lpdiblcb = -1.647835763e-07 wpdiblcb = 2.220446049e-22 ppdiblcb = -1.665334537e-28   drout = 1.478478000e+00 ldrout = -2.828257447e-7   pscbe1 = 6.876139896e+08 lpscbe1 = 3.345779234e+1   pscbe2 = 2.160022972e-08 lpscbe2 = -3.798272305e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.510363785e+00 lbeta0 = 1.189856830e-7   agidl = 1.490566362e-12 lagidl = -8.164949889e-19   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.471888216e-01 lkt1 = 7.296627166e-9   kt2 = -1.323292858e-02 lkt2 = -1.178601122e-8   at = 3.656378506e+03 lat = 1.912648063e-2   ute = 5.522314189e-01 lute = -4.129603001e-07 pute = 4.440892099e-28   ua1 = 5.118987964e-09 lua1 = -1.436452236e-15   ub1 = -4.874445755e-18 lub1 = 1.401068390e-24   uc1 = -2.896530271e-10 luc1 = 5.710342159e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.124 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.093861981e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.395152963e-9   k1 = -1.146151992e+00 lk1 = 5.133688331e-7   k2 = 6.230107875e-01 lk2 = -1.953272252e-07 pk2 = -1.110223025e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.298339775e+00 ldsub = -4.507565858e-07 wdsub = -7.105427358e-21 pdsub = -1.776356839e-27   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.183911471e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.464803694e-8   nfactor = {3.004916136e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.275863248e-7   eta0 = 1.303176041e+00 leta0 = -2.421434955e-7   etab = 8.205958913e-02 letab = -2.445667575e-08 wetab = -3.642919300e-23 petab = 1.019150042e-29   u0 = 6.103225017e-03 lu0 = -2.712861420e-10   ua = -3.514559338e-10 lua = -1.495126584e-16   ub = 8.058113014e-20 lub = 1.468606346e-25   uc = -1.104479542e-12 luc = 3.414877488e-20   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.507369557e+04 lvsat = 5.170207140e-2   a0 = -1.009091321e+00 la0 = 4.835371091e-7   ags = 2.340909297e+00 lags = -2.484818632e-7   a1 = 0.0   a2 = 1.260655052e+00 la2 = -1.383561245e-7   b0 = 0.0   b1 = 0.0   keta = -1.341928945e-01 lketa = 3.051075782e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.867438868e-01 lpclm = -1.475257352e-8   pdiblc1 = 1.128217938e+00 lpdiblc1 = -2.154664579e-07 wpdiblc1 = -3.552713679e-21   pdiblc2 = 2.458828319e-02 lpdiblc2 = -4.767905223e-9   pdiblcb = 2.018475069e-01 lpdiblcb = -1.458702528e-7   drout = -1.004957015e+00 ldrout = 4.566791170e-7   pscbe1 = 7.998864010e+08 lpscbe1 = 2.587504433e-2   pscbe2 = 1.417765344e-08 lpscbe2 = -1.588014653e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.072660264e+01 lbeta0 = -5.409548430e-7   agidl = -1.814317104e-12 lagidl = 1.676166850e-19   bgidl = 2.023190692e+09 lbgidl = -2.330572499e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.659790950e-01 lkt1 = -1.688559918e-8   kt2 = 7.708376428e-02 lkt2 = -3.868006443e-8   at = 1.603330687e+05 lat = -2.752792079e-2   ute = -3.278276177e+00 lute = 7.276690992e-7   ua1 = -1.065189355e-09 lua1 = 4.050411654e-16   ub1 = 7.270196065e-19 lub1 = -2.669079585e-25 pub1 = -3.851859889e-46   uc1 = -3.431547777e-10 luc1 = 7.303490536e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.125 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.9e-07 wmax = 8.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.760176856e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.688950441e-07 wvth0 = 5.276667931e-07 pvth0 = -1.291596393e-13   k1 = 2.702788415e-01 lk1 = 2.049772877e-07 wk1 = 6.332768261e-07 pk1 = -1.550103351e-13   k2 = -7.601578035e-02 lk2 = -3.880125559e-08 wk2 = -7.219006315e-08 pk2 = 1.767032271e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.985721427e+00 ldsub = -6.526526730e-07 wdsub = -2.016371197e-06 pdsub = 4.935572598e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {1.021546984e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.047175391e-08 wvoff = -2.486172503e-07 pvoff = 6.085528743e-14   nfactor = {-1.020358112e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.988537674e-06 wnfactor = 9.233083545e-06 pnfactor = -2.260028025e-12   eta0 = 5.967579281e+00 leta0 = -1.401945192e-06 weta0 = -4.331307355e-06 peta0 = 1.060195758e-12   etab = 5.438140020e-01 letab = -1.393079375e-07 wetab = -4.303919012e-07 petab = 1.053491776e-13   u0 = -5.413085681e-02 lu0 = 1.445226378e-08 wu0 = 4.519489773e-08 pu0 = -1.106258109e-14   ua = -2.826845699e-08 lua = 6.672712390e-15 wua = 2.061533523e-14 pua = -5.046118681e-21   ub = 2.398948524e-17 lub = -5.694480417e-24 wub = -1.759308964e-23 pub = 4.306348516e-30   uc = -2.889493329e-10 luc = 7.049392144e-17 wuc = 2.177908724e-16 puc = -5.330976079e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.067783473e+06 lvsat = -1.195938755e+00 wvsat = -5.548601792e+00 pvsat = 1.358159004e-6   a0 = -4.309906268e+00 la0 = 1.327582907e-06 wa0 = 4.101565413e-06 pa0 = -1.003960674e-12   ags = 1.250000072e+00 lags = -1.545609507e-14   a1 = 0.0   a2 = 2.874371777e+00 la2 = -5.436798531e-07 wa2 = -1.679698100e-06 pa2 = 4.111481025e-13   b0 = 0.0   b1 = 0.0   keta = -2.824694216e-01 lketa = 6.908231687e-08 wketa = 2.134298363e-07 pketa = -5.224228818e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.939684161e-01 lpclm = 6.855483163e-09 wpclm = 2.117994041e-08 ppclm = -5.184319915e-15   pdiblc1 = 4.203168758e+00 lpdiblc1 = -9.842188961e-07 wpdiblc1 = -3.040742876e-06 ppdiblc1 = 7.442978374e-13   pdiblc2 = -5.261860444e-02 lpdiblc2 = 1.377455782e-08 wpdiblc2 = 4.255646371e-08 ppdiblc2 = -1.041675840e-14   pdiblcb = -1.673698382e+01 lpdiblcb = 3.989445150e-06 wpdiblcb = 1.232538432e-05 ppdiblcb = -3.016945946e-12   drout = 1.000001179e+00 ldrout = -2.533148233e-13   pscbe1 = 8.000000009e+08 lpscbe1 = -1.950988770e-7   pscbe2 = -4.052016629e-08 lpscbe2 = 1.168212261e-14 wpscbe2 = 3.609189844e-14 ppscbe2 = -8.834394441e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.405059949e+00 lbeta0 = -1.307342537e-08 wbeta0 = -4.039236401e-08 pbeta0 = 9.887040900e-15   agidl = -2.354088249e-10 lagidl = 5.735822241e-17 wagidl = 1.772081432e-16 pagidl = -4.337612325e-23   bgidl = 1.000000355e+09 lbgidl = -7.620811462e-5   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.607614644e+00 lkt1 = 2.612979846e-07 wkt1 = 8.072797045e-07 pkt1 = -1.976018897e-13   kt2 = 8.832508118e-01 lkt2 = -2.388964923e-07 wkt2 = -7.380703883e-07 pkt2 = 1.806611793e-13   at = -4.537194784e+05 lat = 1.207222435e-01 wat = 3.729712017e-01 pat = -9.129402589e-8   ute = -9.382409569e+00 lute = 2.276117975e-06 wute = 7.032062890e-06 pute = -1.721273194e-12   ua1 = -7.734750384e-09 lua1 = 2.067813237e-15 wua1 = 6.388505373e-15 pua1 = -1.563746403e-21   ub1 = 7.254612413e-18 lub1 = -1.884620178e-24 wub1 = -5.822531841e-24 pub1 = 1.425210231e-30   uc1 = -1.805199625e-10 luc1 = 3.867693277e-17 wuc1 = 1.194923185e-16 puc1 = -2.924873226e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.126 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.127 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.143767018e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.319531148e-7   k1 = 4.210177391e-01 lk1 = 2.132656424e-7   k2 = 5.626381206e-02 lk2 = -3.000267020e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 6.776263578e-27 pcit = 4.743384505e-32   voff = {-1.699412101e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.680610028e-7   nfactor = {1.682760886e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.726492433e-7   eta0 = 0.08   etab = -0.07   u0 = 6.320637964e-03 lu0 = 3.088464059e-8   ua = -7.269192156e-10 lua = 1.507603820e-16   ub = 1.320154755e-19 lub = 9.547120828e-24   uc = -1.283886196e-10 luc = 4.555983095e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.640088689e+04 lvsat = 1.077670413e+0   a0 = 1.632011387e+00 la0 = -3.368254479e-6   ags = 2.730837312e-04 lags = 2.265737709e-6   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 4.581250717e-08 lb0 = -3.686887499e-13   b1 = -6.681756343e-09 lb1 = 5.377327165e-14   keta = 4.028268441e-02 lketa = -3.392369294e-07 wketa = 5.551115123e-23   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 ppclm = 1.332267630e-27   pdiblc1 = 0.39   pdiblc2 = 1.919546137e-03 lpdiblc2 = -1.287843679e-8   pdiblcb = -2.718651916e-01 lpdiblcb = 9.395428170e-7   drout = 0.56   pscbe1 = 8.000326941e+08 lpscbe1 = -6.554436787e-1   pscbe2 = 1.316918687e-08 lpscbe2 = -6.231974900e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.590871467e+01 lbeta0 = -3.189343322e-4   agidl = 2.876157201e-09 lagidl = -1.956461964e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = -4.267601714e-01 legidl = 1.056036940e-05 pegidl = -1.421085472e-26   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.365589613e-01 lkt1 = -3.390156381e-8   kt2 = -6.269565276e-02 lkt2 = 8.319130491e-8   at = 1.185992956e+05 lat = -9.544604462e-1   ute = -4.992636630e-02 lute = -6.626518113e-7   ua1 = 2.269582021e-09 lua1 = -3.596210395e-15   ub1 = -1.572949839e-18 lub1 = 6.897433758e-24   uc1 = -4.389120218e-11 luc1 = 2.827177762e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.128 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.116193739e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004956719e-8   k1 = 4.557220442e-01 lk1 = -6.602679656e-8   k2 = 1.651207896e-02 lk2 = 1.988630180e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.945126661e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.031545343e-8   nfactor = {2.170281296e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.250805327e-6   eta0 = 0.08   etab = -0.07   u0 = 1.011539359e-02 lu0 = 3.453011740e-10   ua = -7.344378443e-10 lua = 2.112686142e-16   ub = 1.372629945e-18 lub = -4.370652867e-25   uc = -7.083236070e-11 luc = -7.601512165e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.684584524e+05 lvsat = -8.703544119e-1   a0 = 1.311480996e+00 la0 = -7.886980138e-7   ags = 2.600278215e-01 lags = 1.752900236e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = -8.302254081e-04 lketa = -8.369481521e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.413146246e-01 lpclm = -8.076396481e-7   pdiblc1 = 0.39   pdiblc2 = -1.408020623e-03 lpdiblc2 = 1.390107179e-08 ppdiblc2 = 1.387778781e-29   pdiblcb = -2.499697493e-01 lpdiblcb = 7.633332238e-7   drout = 0.56   pscbe1 = 1.229788221e+09 lpscbe1 = -3.459231233e+3   pscbe2 = -1.725188617e-08 lpscbe2 = 1.825022021e-13 ppscbe2 = 1.058791184e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.412401616e+00 lbeta0 = 2.306643359e-5   agidl = 6.934301025e-10 lagidl = -1.998523059e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 1.680280514e+00 legidl = -6.396619959e-6   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.059014363e-01 lkt1 = -2.806264270e-7   kt2 = -4.836885543e-02 lkt2 = -3.210753648e-8   at = -9.175901148e+04 lat = 7.384558786e-1   ute = -1.649176185e-01 lute = 2.627719131e-07 wute = -4.440892099e-22   ua1 = 5.627777271e-10 lua1 = 1.013976653e-14   ub1 = 8.332058653e-19 lub1 = -1.246676596e-23 pub1 = -1.232595164e-44   uc1 = -1.166592640e-11 luc1 = 2.337600749e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.129 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.111039678e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081291238e-8   k1 = 4.428479747e-01 lk1 = -1.391545980e-8   k2 = 2.073291406e-02 lk2 = 2.801311033e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.658362304e-01 ldsub = -1.237956247e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.236655549e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.768888085e-8   nfactor = {7.189959202e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.623671336e-6   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411614599e-01 letab = 2.880455783e-7   u0 = 9.794114274e-03 lu0 = 1.645767538e-9   ua = -8.034943736e-10 lua = 4.907939071e-16   ub = 1.317951877e-18 lub = -2.157407696e-25   uc = -7.563850438e-11 luc = 1.185267607e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 53438.0   a0 = 1.119075365e+00 la0 = -9.883308607e-9   ags = 1.669094080e-01 lags = 5.522124099e-7   a1 = 0.0   a2 = 0.8   b0 = 0.0   b1 = 0.0   keta = 6.691932714e-03 lketa = -3.881748511e-08 pketa = -2.775557562e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.631374861e-01 lpclm = 2.448601494e-06 wpclm = -2.220446049e-22   pdiblc1 = 0.39   pdiblc2 = 3.660588932e-03 lpdiblc2 = -6.615519251e-9   pdiblcb = -9.864685163e-02 lpdiblcb = 1.508121816e-7   drout = 0.56   pscbe1 = -5.182772163e+07 lpscbe1 = 1.728461741e+3   pscbe2 = 4.676025648e-08 lpscbe2 = -7.660454858e-14 ppscbe2 = -2.117582368e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.150191084e+01 lbeta0 = -9.678079613e-6   agidl = 2.707512342e-10 lagidl = -2.876141029e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.816907301e-01 lkt1 = 2.615158188e-8   kt2 = -6.033409286e-02 lkt2 = 1.632505246e-8   at = 1.024343241e+05 lat = -4.759505013e-2   ute = -1.331299278e-01 lute = 1.341024937e-7   ua1 = 3.326741149e-09 lua1 = -1.048135508e-15   ub1 = -2.849462571e-18 lub1 = 2.439847267e-24   uc1 = 1.847362934e-11 luc1 = -9.862213274e-17 puc1 = -5.169878828e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.130 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124641429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.704041437e-8   k1 = 3.520889946e-01 lk1 = 1.719385105e-7   k2 = 5.600423158e-02 lk2 = -6.942641121e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.788075222e-01 ldsub = 1.106016613e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.001369456e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.924169099e-10   nfactor = {2.364174723e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.452846867e-7   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = 1.734723476e-24 peta0 = -1.387778781e-28   etab = 8.643192988e-01 letab = -1.770952782e-06 wetab = 7.580741590e-22 petab = 7.754213938e-28   u0 = 1.144702164e-02 lu0 = -1.739014839e-9   ua = -4.031024632e-11 lua = -1.072035469e-15   ub = 5.421819995e-19 lub = 1.372861392e-24   uc = -7.521595276e-11 luc = 1.098738541e-17 wuc = 2.067951531e-31   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.978542095e+04 lvsat = -1.299808994e-2   a0 = 1.428287075e+00 la0 = -6.430793195e-7   ags = 1.532493533e-01 lags = 5.801851283e-7   a1 = 0.0   a2 = 5.904554777e-01 la2 = 4.291000341e-7   b0 = 0.0   b1 = 0.0   keta = -1.076463397e-02 lketa = -3.070364262e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.508138941e-01 lpclm = 3.722572068e-7   pdiblc1 = 7.577690250e-01 lpdiblc1 = -7.531082152e-7   pdiblc2 = 0.00043   pdiblcb = -0.025   drout = 9.897900000e-02 ldrout = 9.440672783e-7   pscbe1 = 7.984623780e+08 lpscbe1 = -1.274106762e+1   pscbe2 = 9.534760526e-09 lpscbe2 = -3.751086118e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 5.840666904e+00 lbeta0 = 1.914874189e-6   agidl = -2.655058546e-10 lagidl = 8.105197571e-16 pagidl = 4.135903063e-37   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.582905950e-01 lkt1 = -2.176662973e-8   kt2 = -5.634649868e-02 lkt2 = 8.159356780e-9   at = 9.745498753e+04 lat = -3.739848929e-2   ute = 9.597179901e-01 lute = -2.103804152e-06 wute = 6.661338148e-22 pute = -8.881784197e-28   ua1 = 6.215248388e-09 lua1 = -6.963148420e-15   ub1 = -4.332849657e-18 lub1 = 5.477490257e-24   uc1 = -1.309081232e-10 luc1 = 2.072780856e-16 wuc1 = 1.033975766e-31   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.131 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140123256e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.326188593e-8   k1 = 5.232439484e-01 lk1 = -7.393371107e-9   k2 = -1.226088730e-02 lk2 = 2.100073728e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.277500803e+00 ldsub = -5.246443427e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.926698888e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.316212391e-9   nfactor = {1.185783805e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.894038578e-7   eta0 = -3.486985538e-02 leta0 = 2.670462627e-7   etab = -1.729964684e+00 letab = 9.472731180e-7   u0 = 1.389723133e-02 lu0 = -4.306283297e-9   ua = -9.132162872e-10 lua = -1.574263421e-16   ub = 2.527606944e-18 lub = -7.074172299e-25   uc = -1.014940739e-10 luc = 3.852094380e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.311994564e+04 lvsat = 1.157790805e-1   a0 = 8.881460474e-01 la0 = -7.713305401e-8   ags = 1.120744391e-01 lags = 6.233271741e-7   a1 = 0.0   a2 = 1.053132798e+00 la2 = -5.568169504e-8   b0 = -9.608784530e-17 lb0 = 1.006784421e-22   b1 = -3.994811609e-20 lb1 = 4.185663734e-26   keta = 1.311717861e-02 lketa = -2.809313044e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.624337286e+00 lpclm = -8.573312648e-07 wpclm = 3.552713679e-21   pdiblc1 = 6.467424655e-02 lpdiblc1 = -2.690083368e-8   pdiblc2 = 7.922616047e-04 lpdiblc2 = -3.795686529e-10   pdiblcb = -1.354002314e-02 lpdiblcb = -1.200747726e-8   drout = 1.041454917e+00 ldrout = -4.343542515e-8   pscbe1 = 8.275046100e+08 lpscbe1 = -4.317079225e+1   pscbe2 = 3.162763138e-09 lpscbe2 = 6.301310952e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 6.507657499e+00 lbeta0 = 1.216018119e-6   agidl = 1.064658721e-09 lagidl = -5.831934307e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.190246567e-01 lkt1 = -6.290849829e-8   kt2 = -6.368883441e-02 lkt2 = 1.585247260e-8   at = 8.716611382e+04 lat = -2.661806463e-02 wat = 2.328306437e-16   ute = -1.975547800e+00 lute = 9.716939615e-07 wute = -3.552713679e-21   ua1 = -3.637135874e-09 lua1 = 3.359933500e-15   ub1 = 4.413339682e-18 lub1 = -3.686548278e-24 pub1 = 1.540743956e-45   uc1 = 3.433541843e-10 luc1 = -2.896421036e-16 wuc1 = -2.067951531e-31   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.132 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.083758130e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.386478892e-9   k1 = 4.286126363e-01 lk1 = 4.444329585e-8   k2 = 2.077621672e-02 lk2 = -1.599682593e-08 pk2 = 1.387778781e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.339715233e-01 ldsub = 3.033024110e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.158159998e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.362648555e-9   nfactor = {1.886976015e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.053082948e-7   eta0 = 4.081427101e-01 leta0 = 2.437505465e-8   etab = -1.347621329e-03 letab = 3.799063485e-10   u0 = 7.040683625e-03 lu0 = -5.504378792e-10   ua = -1.613983779e-09 lua = 2.264365708e-16   ub = 2.025147933e-18 lub = -4.321827452e-25   uc = -6.712093967e-11 luc = 1.969220019e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.716932025e+05 lvsat = -1.284569167e-2   a0 = 9.052648244e-01 la0 = -8.651029208e-8   ags = 9.445453886e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.136650759e+00 la2 = -1.014307462e-7   b0 = 1.921756906e-16 lb0 = -5.722511627e-23   b1 = 7.989623218e-20 lb1 = -2.379110054e-26   keta = -4.583734636e-02 lketa = 4.200684472e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.292099820e-01 lpclm = 3.771055897e-07 ppclm = -3.330669074e-28   pdiblc1 = -4.478501477e-01 lpdiblc1 = 2.538472164e-07 wpdiblc1 = -2.775557562e-22 ppdiblc1 = -5.551115123e-29   pdiblc2 = -9.997833428e-03 lpdiblc2 = 5.530975654e-09 wpdiblc2 = 8.673617380e-25 ppdiblc2 = -6.179952383e-30   pdiblcb = 2.653629919e-01 lpdiblcb = -1.647835763e-07 ppdiblcb = -5.551115123e-29   drout = 1.478478000e+00 ldrout = -2.828257447e-7   pscbe1 = 6.876139896e+08 lpscbe1 = 3.345779234e+1   pscbe2 = 2.160022972e-08 lpscbe2 = -3.798272305e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.510363785e+00 lbeta0 = 1.189856830e-7   agidl = 1.490566362e-12 lagidl = -8.164949889e-19   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.471888216e-01 lkt1 = 7.296627166e-9   kt2 = -1.323292858e-02 lkt2 = -1.178601122e-8   at = 3.656378506e+03 lat = 1.912648063e-2   ute = 5.522314189e-01 lute = -4.129603001e-07 pute = -2.220446049e-28   ua1 = 5.118987964e-09 lua1 = -1.436452236e-15   ub1 = -4.874445755e-18 lub1 = 1.401068390e-24   uc1 = -2.896530271e-10 luc1 = 5.710342159e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.133 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.093861981e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.395152963e-9   k1 = -1.146151992e+00 lk1 = 5.133688331e-7   k2 = 6.230107875e-01 lk2 = -1.953272252e-07 pk2 = -1.110223025e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.298339775e+00 ldsub = -4.507565858e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.183911471e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.464803694e-8   nfactor = {3.004916136e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.275863248e-7   eta0 = 1.303176041e+00 leta0 = -2.421434955e-7   etab = 8.205958913e-02 letab = -2.445667575e-08 wetab = -6.158268340e-23 petab = -2.775557562e-29   u0 = 6.103225017e-03 lu0 = -2.712861420e-10   ua = -3.514559338e-10 lua = -1.495126584e-16   ub = 8.058113014e-20 lub = 1.468606346e-25   uc = -1.104479542e-12 luc = 3.414877488e-20   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.507369557e+04 lvsat = 5.170207140e-2   a0 = -1.009091321e+00 la0 = 4.835371091e-7   ags = 2.340909297e+00 lags = -2.484818632e-7   a1 = 0.0   a2 = 1.260655052e+00 la2 = -1.383561245e-7   b0 = 0.0   b1 = 0.0   keta = -1.341928945e-01 lketa = 3.051075782e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.867438868e-01 lpclm = -1.475257352e-8   pdiblc1 = 1.128217938e+00 lpdiblc1 = -2.154664579e-7   pdiblc2 = 2.458828319e-02 lpdiblc2 = -4.767905223e-9   pdiblcb = 2.018475069e-01 lpdiblcb = -1.458702528e-7   drout = -1.004957015e+00 ldrout = 4.566791170e-7   pscbe1 = 7.998864010e+08 lpscbe1 = 2.587504434e-2   pscbe2 = 1.417765344e-08 lpscbe2 = -1.588014653e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.072660264e+01 lbeta0 = -5.409548430e-7   agidl = -1.814317104e-12 lagidl = 1.676166850e-19   bgidl = 2.023190692e+09 lbgidl = -2.330572499e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.659790950e-01 lkt1 = -1.688559918e-8   kt2 = 7.708376428e-02 lkt2 = -3.868006443e-8   at = 1.603330687e+05 lat = -2.752792079e-2   ute = -3.278276177e+00 lute = 7.276690992e-7   ua1 = -1.065189355e-09 lua1 = 4.050411654e-16 pua1 = 4.135903063e-37   ub1 = 7.270196065e-19 lub1 = -2.669079585e-25   uc1 = -3.431547777e-10 luc1 = 7.303490536e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.134 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.5e-07 wmax = 7.9e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.024322225e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.122377318e-08 wvth0 = -6.734387086e-09 pvth0 = 1.648409599e-15   k1 = 2.752502636e-01 lk1 = 2.037604078e-07 wk1 = 6.296664203e-07 pk1 = -1.541265980e-13   k2 = 7.135804066e-02 lk2 = -7.487468263e-08 wk2 = -1.792176479e-07 pk2 = 4.386799977e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.969892279e+00 ldsub = -6.487780933e-07 wdsub = -2.004875564e-06 pdsub = 4.907434161e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {1.021532160e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.047139106e-08 wvoff = -2.486161737e-07 pvoff = 6.085502392e-14   nfactor = {-1.020358191e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.988537867e-06 wnfactor = 9.233084117e-06 pnfactor = -2.260028165e-12   eta0 = 5.967580365e+00 leta0 = -1.401945457e-06 weta0 = -4.331308143e-06 peta0 = 1.060195951e-12   etab = 5.404352903e-01 letab = -1.384809134e-07 wetab = -4.279381726e-07 petab = 1.047485662e-13   u0 = -4.021109693e-02 lu0 = 1.104505456e-08 wu0 = 3.508592266e-08 pu0 = -8.588156720e-15   ua = -2.826858426e-08 lua = 6.672743542e-15 wua = 2.061542766e-14 pua = -5.046141305e-21   ub = 2.399089283e-17 lub = -5.694824959e-24 wub = -1.759411187e-23 pub = 4.306598734e-30   uc = -2.872396061e-10 luc = 7.007542307e-17 wuc = 2.165492141e-16 puc = -5.300583387e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.972765371e+07 lvsat = 1.221661438e+01 wvsat = 3.424559814e+01 pvsat = -8.382466285e-6   a0 = -4.309907218e+00 la0 = 1.327583140e-06 wa0 = 4.101566102e-06 pa0 = -1.003960843e-12   ags = 1.250000072e+00 lags = -1.545608797e-14   a1 = 0.0   a2 = 2.861185619e+00 la2 = -5.404522113e-07 wa2 = -1.670121890e-06 pa2 = 4.088040857e-13   b0 = 0.0   b1 = 0.0   keta = -2.824694192e-01 lketa = 6.908231629e-08 wketa = 2.134298346e-07 pketa = -5.224228776e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.941346852e-01 lpclm = 6.814784623e-09 wpclm = 2.105919041e-08 ppclm = -5.154763332e-15   pdiblc1 = 4.179297971e+00 lpdiblc1 = -9.783759242e-07 wpdiblc1 = -3.023407146e-06 ppdiblc1 = 7.400544842e-13   pdiblc2 = -5.228452282e-02 lpdiblc2 = 1.369278299e-08 wpdiblc2 = 4.231384295e-08 ppdiblc2 = -1.035737091e-14   pdiblcb = -1.664022568e+01 lpdiblcb = 3.965761177e-06 wpdiblcb = 1.225511546e-05 ppdiblcb = -2.999745886e-12   drout = 1.000001179e+00 ldrout = -2.533148518e-13 wdrout = -8.526512829e-20 pdrout = 2.131628207e-26   pscbe1 = 8.000000009e+08 lpscbe1 = -1.950988770e-7   pscbe2 = -4.023683355e-08 lpscbe2 = 1.161276984e-14 wpscbe2 = 3.588613314e-14 ppscbe2 = -8.784028238e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.404742856e+00 lbeta0 = -1.299580899e-08 wbeta0 = -4.016208110e-08 pbeta0 = 9.830673402e-15   agidl = -1.327055042e-10 lagidl = 3.221901709e-17 wagidl = 1.026217052e-16 pagidl = -2.511922789e-23   bgidl = 1.000000355e+09 lbgidl = -7.620812225e-5   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.607616049e+00 lkt1 = 2.612983287e-07 wkt1 = 8.072807254e-07 pkt1 = -1.976021396e-13   kt2 = 8.774567273e-01 lkt2 = -2.374782453e-07 wkt2 = -7.338625387e-07 pkt2 = 1.796312029e-13   at = -4.507915372e+05 lat = 1.200055567e-01 wat = 3.708448371e-01 pat = -9.077354500e-8   ute = -9.327205665e+00 lute = 2.262605439e-06 wute = 6.991972048e-06 pute = -1.711459958e-12   ua1 = -7.684598609e-09 lua1 = 2.055537336e-15 wua1 = 6.352083549e-15 pua1 = -1.554831251e-21   ub1 = 7.208903708e-18 lub1 = -1.873431830e-24 wub1 = -5.789336717e-24 pub1 = 1.417084895e-30   uc1 = -1.795819103e-10 luc1 = 3.844732103e-17 wuc1 = 1.188110749e-16 puc1 = -2.908198087e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.135 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.136 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.391472862e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.197904136e-06 wvth0 = 1.699836765e-07 pvth0 = -3.407794501e-12   k1 = 4.721684590e-01 lk1 = -8.121924824e-07 wk1 = -3.510126086e-08 pk1 = 7.037021799e-13   k2 = 3.575905468e-02 lk2 = 1.110480602e-07 wk2 = 1.407102066e-08 pk2 = -2.820926562e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = -2.541098842e-27 pcit = 1.355252716e-32   voff = {-3.671690496e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.685918348e-06 wvoff = 1.353440548e-07 pvoff = -2.713347158e-12   nfactor = {6.075466187e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.319026507e-05 wnfactor = 1.113072575e-06 pnfactor = -2.231462855e-11   eta0 = 0.08   etab = -0.07   u0 = 9.347517593e-03 lu0 = -2.979756116e-08 wu0 = -2.077141662e-09 pu0 = 4.164206867e-14   ua = -1.557939953e-09 lua = 1.681087714e-14 wua = 5.702730225e-16 pua = -1.143270524e-20   ub = 1.218603947e-18 lub = -1.223656037e-23 wub = -7.456517802e-25 pub = 1.494865912e-29   uc = -4.304485922e-10 luc = 6.511228675e-15 wuc = 2.072832191e-16 puc = -4.155567337e-21   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -8.205399596e+05 lvsat = 1.805694994e+01 wvsat = 5.811979110e-01 pvsat = -1.165172495e-5   a0 = 1.695517019e+00 la0 = -4.641401100e-06 wa0 = -4.357959684e-08 pa0 = 8.736739521e-13   ags = -1.430854157e+00 lags = 3.095665463e-05 wags = 9.820853088e-07 pags = -1.968862530e-11   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = -9.627917961e-07 lb0 = 1.985158339e-11 wb0 = 6.921365482e-13 pb0 = -1.387579779e-17   b1 = -5.119311450e-09 lb1 = 2.244972799e-14 wb1 = -1.072199684e-15 pb1 = 2.149521801e-20   keta = 1.170910408e-01 lketa = -1.879073577e-06 wketa = -5.270835204e-08 pketa = 1.056685182e-12   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 ppclm = -6.661338148e-28   pdiblc1 = 0.39   pdiblc2 = 2.021311486e-03 lpdiblc2 = -1.491860562e-08 wpdiblc2 = -6.983463934e-11 ppdiblc2 = 1.400029137e-15   pdiblcb = -8.682078835e-01 lpdiblcb = 1.289488693e-05 wpdiblcb = 4.092294382e-07 ppdiblcb = -8.204139700e-12   drout = 0.56   pscbe1 = 8.004487146e+08 lpscbe1 = -8.995728530e+00 wpscbe1 = -2.854865617e-01 ppscbe1 = 5.723370354e-6   pscbe2 = 6.803838913e-08 lpscbe2 = -1.162325170e-12 wpscbe2 = -3.765300241e-14 ppscbe2 = 7.548589203e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 1.793004239e+01 lbeta0 = 2.419757945e-04 wbeta0 = 1.919986024e-05 pbeta0 = -3.849144780e-10   agidl = 3.658102371e-09 lagidl = -3.524088047e-14 wagidl = -5.365957979e-16 pagidl = 1.075755182e-20   bgidl = 1000000000.0   cgidl = 300.0   egidl = -7.129593719e+00 legidl = 1.449372682e-04 wegidl = 4.599698871e-06 pegidl = -9.221372803e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.366563594e-01 lkt1 = -2.036726448e-06 wkt1 = -6.855636228e-08 pkt1 = 1.374402526e-12   kt2 = -3.027344063e-02 lkt2 = -5.668019089e-07 wkt2 = -2.224915948e-08 pkt2 = 4.460461431e-13   at = 6.456587741e+05 lat = -1.152083028e+01 wat = -3.616850801e-01 pat = 7.250981106e-6   ute = -7.865937086e+00 lute = 1.560309725e-04 wute = 5.363596668e-06 pute = -1.075281792e-10   ua1 = -1.695805897e-08 lua1 = 3.818752100e-13 wua1 = 1.319462253e-14 pua1 = -2.645228238e-19   ub1 = 1.217300178e-17 lub1 = -2.686783114e-22 wub1 = -9.432911871e-24 pub1 = 1.891088948e-28   uc1 = 6.019437063e-10 luc1 = -1.266483516e-14 wuc1 = -4.431925809e-16 puc1 = 8.885025144e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.137 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-8.023312090e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.566246731e-07 wvth0 = -2.153825114e-07 pvth0 = -3.064541281e-13   k1 = 3.955361438e-01 lk1 = -1.954728512e-07 wk1 = 4.130149082e-08 pk1 = 8.883002496e-14   k2 = 5.377679140e-02 lk2 = -3.395463092e-08 wk2 = -2.557223815e-08 pk2 = 3.694737094e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {4.027421796e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.510153995e-06 wvoff = -4.098553873e-07 pvoff = 1.674295282e-12   nfactor = {1.712703613e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.041553282e-04 wnfactor = -1.026380378e-05 pnfactor = 6.924391257e-11   eta0 = 0.08   etab = -0.07   u0 = 1.785951368e-02 lu0 = -9.830019047e-08 wu0 = -5.314263021e-09 pu0 = 6.769369302e-14   ua = 2.321959749e-09 lua = -1.441368268e-14 wua = -2.097397833e-15 pua = 1.003610958e-20   ub = 1.043683610e-19 lub = -3.269443077e-24 wub = 8.703216835e-25 pub = 1.943668276e-30   uc = 3.894654781e-10 luc = -8.725528187e-17 wuc = -3.158711065e-16 puc = 5.466096570e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 2.877049213e+06 lvsat = -1.170041576e+01 wvsat = -1.790098455e+00 pvsat = 7.431934662e-6   a0 = 3.125886013e+00 la0 = -1.615268893e-05 wa0 = -1.245102784e-06 pa0 = 1.054326222e-11   ags = 3.004452091e+00 lags = -4.737692108e-06 wags = -1.883311755e-06 pags = 3.371445554e-12   a1 = 0.0   a2 = 0.8   b0 = 1.120588227e-06 lb0 = 3.085009724e-12 wb0 = -7.689834999e-13 pb0 = -2.117032393e-18   b1 = -4.550106917e-08 lb1 = 3.474330283e-13 wb1 = 3.122428970e-14 pb1 = -2.384196618e-19   keta = -1.073748816e-01 lketa = -7.262233761e-08 wketa = 7.311435254e-08 pketa = 4.409236594e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 8.583273543e+00 lpclm = -6.794184808e-05 wpclm = -5.724519152e-06 ppclm = 4.606964212e-11   pdiblc1 = 0.39   pdiblc2 = -2.226735725e-02 lpdiblc2 = 1.805511354e-07 wpdiblc2 = 1.431434429e-08 ppdiblc2 = -1.143606064e-13   pdiblcb = -5.677008203e-01 lpdiblcb = 1.047647370e-05 wpdiblcb = 2.180372283e-07 ppdiblcb = -6.665467813e-12   drout = 0.56   pscbe1 = 6.698688616e+09 lpscbe1 = -4.747670335e+04 wpscbe1 = -3.752934455e+03 ppscbe1 = 3.020619792e-2   pscbe2 = -4.232129785e-07 lpscbe2 = 2.791155305e-12 wpscbe2 = 2.785834923e-13 ppscbe2 = -1.790141236e-18   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.187661992e-09 lalpha0 = 1.036281399e-14 walpha0 = 8.836348640e-16 palpha0 = -7.111294568e-21   alpha1 = -1.187661992e-09 lalpha1 = 1.036281399e-14 walpha1 = 8.836348640e-16 palpha1 = -7.111294568e-21   beta0 = 3.563288015e+02 lbeta0 = -2.481381279e-03 wbeta0 = -2.421825269e-04 pbeta0 = 1.718632163e-9   agidl = 6.659902202e-10 lagidl = -1.116103510e-14 wagidl = 1.883012533e-17 pagidl = 6.287608963e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 2.178878116e+01 legidl = -8.779130615e-05 wegidl = -1.379909661e-05 pegidl = 5.585563829e-11   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.066915568e-01 lkt1 = -2.277876437e-06 wkt1 = -6.808099404e-08 pkt1 = 1.370576869e-12   kt2 = -1.745435035e-01 lkt2 = 5.942510967e-07 wkt2 = 8.658508113e-08 pkt2 = -4.298273375e-13   at = -1.540127989e+06 lat = 6.069889786e+00 wat = 9.939171403e-01 pat = -3.658600553e-6   ute = 2.221461262e+01 lute = -8.605052342e-05 wute = -1.535754979e-05 pute = 5.923094528e-11   ua1 = 4.565751708e-08 lua1 = -1.220408575e-13 wua1 = -3.094545317e-14 pua1 = 9.070657400e-20   ub1 = -2.601116324e-17 lub1 = 3.861925722e-23 wub1 = 1.842146510e-23 pub1 = -3.505686386e-29   uc1 = -7.257545625e-09 luc1 = 5.058656659e-14 wuc1 = 4.972354517e-15 puc1 = -3.469807940e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.138 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-6.734446492e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.507912147e-08 wvth0 = -3.002917114e-07 pvth0 = 3.723920920e-14   k1 = 1.183952155e+00 lk1 = -3.386803472e-06 wk1 = -5.085694040e-07 pk1 = 2.314583686e-12   k2 = -2.535353885e-01 lk2 = 1.209975928e-06 wk2 = 1.882116858e-07 pk2 = -8.284018519e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.489123398e-01 ldsub = -1.169452146e-06 wdsub = 1.161371531e-08 pdsub = -4.700970647e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-3.204368576e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.171120321e-07 wvoff = 6.640756460e-08 pvoff = -2.535099879e-13   nfactor = {-1.833267270e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.937759465e-05 wnfactor = 1.307386466e-05 pnfactor = -2.522171830e-11   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411777301e-01 letab = 2.881114366e-07 wetab = 1.116516329e-11 petab = -4.519406884e-17   u0 = -2.759200612e-02 lu0 = 8.567733510e-08 wu0 = 2.565555217e-08 pu0 = -5.766515067e-14   ua = -7.103796988e-09 lua = 2.373965979e-14 wua = 4.323469264e-15 pua = -1.595411574e-20   ub = 3.695526850e-18 lub = -1.780564463e-23 wub = -1.631568029e-24 pub = 1.207075491e-29   uc = 6.685958989e-10 luc = -1.217112421e-15 wuc = -5.107174631e-16 puc = 8.433551764e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -3.378889433e+05 lvsat = 1.312930533e+00 wvsat = 2.685410709e-01 pvsat = -9.009749452e-7   a0 = -2.484914548e+00 la0 = 6.558569307e-06 wa0 = 2.473173206e-06 pa0 = -4.507482375e-12   ags = 2.889418240e+00 lags = -4.272060961e-06 wags = -1.868272681e-06 pags = 3.310570764e-12   a1 = 0.0   a2 = 0.8   b0 = 2.493779067e-06 lb0 = -2.473357829e-12 wb0 = -1.711310997e-12 pb0 = 1.697297290e-18   b1 = 3.878031270e-08 lb1 = 6.280957728e-15 wb1 = -2.661229155e-14 pb1 = -4.310194184e-21   keta = -2.008704513e-01 lketa = 3.058266920e-07 wketa = 1.424359499e-07 pketa = -2.365058629e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -1.542711067e+01 lpclm = 2.924678486e-05 wpclm = 1.020013404e-05 ppclm = -1.838977097e-11   pdiblc1 = 0.39   pdiblc2 = 4.491620165e-02 lpdiblc2 = -9.139279471e-08 wpdiblc2 = -2.831092162e-08 ppdiblc2 = 5.817687929e-14   pdiblcb = 4.114871442e+00 lpdiblcb = -8.477525242e-06 wpdiblcb = -2.891451086e-06 ppdiblcb = 5.921041247e-12   drout = 0.56   pscbe1 = -1.089102882e+10 lpscbe1 = 2.372251515e+04 wpscbe1 = 7.438206649e+03 ppscbe1 = -1.509302326e-2   pscbe2 = 5.309623611e-07 lpscbe2 = -1.071131780e-12 wpscbe2 = -3.322749787e-13 ppscbe2 = 6.824764113e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.675323984e-09 lalpha0 = -5.273684071e-15 walpha0 = -1.767269728e-15 palpha0 = 3.618970767e-21   alpha1 = 2.675323984e-09 lalpha1 = -5.273684071e-15 walpha1 = -1.767269728e-15 palpha1 = 3.618970767e-21   beta0 = -5.421957297e+02 lbeta0 = 1.155643855e-03 wbeta0 = 3.799650393e-04 pbeta0 = -7.996812020e-10   agidl = 4.720255204e-09 lagidl = -2.757178755e-14 wagidl = -3.053392009e-15 pagidl = 1.872327291e-20   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.070417073e+00 lkt1 = 8.135126137e-07 wkt1 = 4.040028557e-07 pkt1 = -5.403123356e-13   kt2 = -2.301205697e-02 lkt2 = -1.911410450e-08 wkt2 = -2.561157533e-08 pkt2 = 2.431948356e-14   at = -6.732542753e+05 lat = 2.560980039e+00 wat = 5.323023389e-01 pat = -1.790087700e-6   ute = -6.762002730e-01 lute = 6.606336743e-06 wute = 3.726722491e-07 pute = -4.441454254e-12   ua1 = 8.801259739e-09 lua1 = 2.714497953e-14 wua1 = -3.756789841e-15 pua1 = -1.934701772e-20   ub1 = -1.475136867e-17 lub1 = -6.957857748e-24 wub1 = 8.167468827e-24 pub1 = 6.449005907e-30   uc1 = 1.148485766e-08 luc1 = -2.527846485e-14 wuc1 = -7.868599643e-15 puc1 = 1.727921382e-20   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.139 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-7.223859716e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.514169500e-08 wvth0 = -2.760405671e-07 pvth0 = -1.242167801e-14   k1 = -1.612055820e+00 lk1 = 2.338791759e-06 wk1 = 1.347859024e-06 pk1 = -1.486964039e-12   k2 = 8.013947456e-01 lk2 = -9.502836272e-07 wk2 = -5.115108232e-07 pk2 = 6.044724090e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -7.134939531e+00 ldsub = 1.517968012e-05 wdsub = 4.704897181e-06 pdsub = -9.657798255e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-8.092076228e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.336303991e-08 wvoff = -8.180995994e-08 pvoff = 5.000615337e-14   nfactor = {5.398394028e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.309361779e-07 wnfactor = 1.251917275e-06 pnfactor = -1.013029996e-12   eta0 = 3.370304500e+00 leta0 = -6.900601410e-06 weta0 = -2.470291855e-06 peta0 = 5.058601903e-12   etab = 1.185887448e+01 letab = -2.428529547e-05 wetab = -7.544815588e-06 petab = 1.545006241e-11   u0 = -8.228471453e-03 lu0 = 4.602517289e-08 wu0 = 1.350195297e-08 pu0 = -3.277731407e-14   ua = 4.332156425e-09 lua = 3.214002943e-16 wua = -3.000526549e-15 pua = -9.562202108e-22   ub = -1.105381056e-17 lub = 1.239767979e-23 wub = 7.957541168e-24 pub = -7.565583178e-30   uc = 5.017539703e-10 luc = -8.754576904e-16 wuc = -3.959352242e-16 puc = 6.083069773e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.304631929e+05 lvsat = -6.700367632e-01 wvsat = -3.916173488e-01 pvsat = 4.508809629e-7   a0 = 6.518919416e+00 la0 = -1.187925679e-05 wa0 = -3.493354812e-06 pa0 = 7.710624536e-12   ags = -9.986256867e-01 lags = 3.689778190e-06 wags = 7.904535125e-07 pags = -2.133902266e-12   a1 = 0.0   a2 = -2.075923132e+00 la2 = 5.889243491e-06 wa2 = 1.829754326e-06 pa2 = -3.746925165e-12   b0 = 8.522179398e-08 lb0 = 2.458825540e-12 wb0 = -5.848192213e-14 pb0 = -1.687324768e-18   b1 = 8.690354907e-08 lb1 = -9.226460263e-14 wb1 = -5.963599629e-14 pb1 = 6.331492279e-20   keta = 7.760375976e-02 lketa = -2.644258356e-07 wketa = -6.064121957e-08 pketa = 1.793504878e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -5.562876073e+00 lpclm = 9.047051866e-06 wpclm = 4.126786493e-06 ppclm = -5.952921688e-12   pdiblc1 = 5.362023718e+00 lpdiblc1 = -1.018158587e-05 wpdiblc1 = -3.159586906e-06 ppdiblc1 = 6.470123077e-12   pdiblc2 = 1.349368697e-04 lpdiblc2 = 3.091597713e-10 wpdiblc2 = 2.024817620e-10 ppdiblc2 = -2.121553282e-16   pdiblcb = -2.691511935e+00 lpdiblcb = 5.460416478e-06 wpdiblcb = 1.829845818e-06 ppdiblcb = -3.747112521e-12   drout = -3.415944104e+00 ldrout = 8.141838937e-06 wdrout = 2.412052711e-06 pdrout = -4.939341241e-12   pscbe1 = 7.788966914e+08 lpscbe1 = -1.748665663e+02 wpscbe1 = 1.342660026e+01 ppscbe1 = 1.112557052e-4   pscbe2 = 6.456026751e-09 lpscbe2 = 2.939178536e-15 wpscbe2 = 2.112725636e-15 ppscbe2 = -2.274369898e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 2.135630311e+01 lbeta0 = 1.616091121e-06 wbeta0 = -1.064732606e-05 pbeta0 = 2.050345029e-13   agidl = -8.758005219e-09 lagidl = 2.865719171e-17 wagidl = 5.827824824e-15 pagidl = 5.365391120e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -8.765086498e-01 lkt1 = 4.164317926e-07 wkt1 = 2.869946122e-07 pkt1 = -3.007057798e-13   kt2 = -1.535852359e-02 lkt2 = -3.478681882e-08 wkt2 = -2.812726012e-08 pkt2 = 2.947103997e-14   at = 9.842687581e+05 lat = -8.332541910e-01 wat = -6.085599874e-01 pat = 5.461416499e-7   ute = 6.319866364e+00 lute = -7.720033614e-06 wute = -3.678305339e-06 pute = 3.854036376e-12   ua1 = 4.561894574e-08 lua1 = -4.824935741e-14 wua1 = -2.704007804e-14 pua1 = 2.833191777e-20   ub1 = -3.863628282e-17 lub1 = 4.195307233e-23 wub1 = 2.354011355e-23 pub1 = -2.503071164e-29   uc1 = -1.830176286e-09 luc1 = 1.987728785e-15 wuc1 = 1.166092190e-15 puc1 = -1.221802244e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.140 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-2.609742713e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.483139493e-07 wvth0 = -6.033001663e-07 pvth0 = 3.304727486e-13   k1 = 7.409867799e-01 lk1 = -1.266674507e-07 wk1 = -1.494220988e-07 pk1 = 8.184969016e-14   k2 = -2.119722276e-01 lk2 = 1.114969532e-07 wk2 = 1.370483125e-07 pk2 = -7.507163936e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.505746038e+01 ldsub = -8.072961702e-06 wdsub = -9.456249223e-06 pdsub = 5.179896918e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-8.858766178e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.532985430e-08 wvoff = -7.142455481e-08 pvoff = 3.912458551e-14   nfactor = {3.152396536e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.662661801e-07 wnfactor = 5.973952538e-07 pnfactor = -3.272381852e-13   eta0 = -7.234452080e+00 leta0 = 4.210797416e-06 weta0 = 4.940583709e-06 peta0 = -2.706328241e-12   etab = -2.371900996e+01 letab = 1.299232239e-05 wetab = 1.508958652e-05 petab = -8.265698253e-12   u0 = 6.819462724e-02 lu0 = -3.404903934e-08 wu0 = -3.726061059e-08 pu0 = 2.041043097e-14   ua = 1.103637777e-08 lua = -6.703115228e-15 wua = -8.200193831e-15 pua = 4.491861176e-21   ub = 2.772615266e-19 lub = 5.252657312e-25 wub = 1.544259037e-24 pub = -8.459064938e-31   uc = -6.653149034e-10 luc = 3.473678987e-16 wuc = 3.869118954e-16 puc = -2.119406635e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.813134871e+05 lvsat = 1.805225477e-01 wvsat = 8.110819037e-02 pvsat = -4.442903898e-8   a0 = -1.091653429e+01 la0 = 6.389175717e-06 wa0 = 8.100749396e-06 pa0 = -4.437388000e-12   ags = 3.917448822e+00 lags = -1.461161779e-06 wags = -2.611369674e-06 pags = 1.430443023e-12   a1 = 0.0   a2 = 6.385890017e+00 la2 = -2.976832781e-06 wa2 = -3.659508652e-06 pa2 = 2.004587352e-12   b0 = 5.096237610e-06 lb0 = -2.791591557e-12 wb0 = -3.497201328e-12 pb0 = 1.915679457e-18   b1 = -2.418472995e-09 lb1 = 1.324779045e-15 wb1 = 1.659633560e-15 pb1 = -9.091057735e-22   keta = -3.244133766e-01 lketa = 1.567976694e-07 wketa = 2.316242680e-07 pketa = -1.268779834e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.371938593e+00 lpclm = -3.457948571e-06 wpclm = -3.257955941e-06 ppclm = 1.784626815e-12   pdiblc1 = -9.143835138e+00 lpdiblc1 = 5.017290395e-06 wpdiblc1 = 6.319173812e-06 ppdiblc1 = -3.461485435e-12   pdiblc2 = 7.922616047e-04 lpdiblc2 = -3.795686529e-10   pdiblcb = 5.319483847e+00 lpdiblcb = -2.933304628e-06 wpdiblcb = -3.659691637e-06 ppdiblcb = 2.004687586e-12   drout = 8.071301124e+00 ldrout = -3.894209432e-06 wdrout = -4.824105423e-06 pdrout = 2.642524348e-12   pscbe1 = 4.622527380e+08 lpscbe1 = 1.569050519e+02 wpscbe1 = 2.506475226e+02 ppscbe1 = -1.372984467e-4   pscbe2 = 3.339696871e-09 lpscbe2 = 6.204391076e-15 wpscbe2 = -1.214175894e-16 ppscbe2 = 6.650952005e-23   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 3.842388281e+01 lbeta0 = -1.626689220e-05 wbeta0 = -2.190193513e-05 pbeta0 = 1.199733251e-11   agidl = -1.829552345e-08 lagidl = 1.002183036e-14 wagidl = 1.328557653e-14 pagidl = -7.277506686e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.190246567e-01 lkt1 = -6.290849829e-8   kt2 = -6.368883441e-02 lkt2 = 1.585247260e-8   at = 3.538173073e+05 lat = -1.726829222e-01 wat = -1.829845818e-01 pat = 1.002343793e-7   ute = -1.975547800e+00 lute = 9.716939615e-7   ua1 = -3.637135874e-09 lua1 = 3.359933500e-15 wua1 = -3.308722450e-30   ub1 = 5.479944456e-18 lub1 = -4.270807708e-24 wub1 = -7.319383273e-25 pub1 = 4.009375173e-31   uc1 = 3.433541843e-10 luc1 = -2.896421036e-16 puc1 = 1.033975766e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.141 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.083758130e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.386478892e-9   k1 = 4.286126363e-01 lk1 = 4.444329585e-8   k2 = 2.077621672e-02 lk2 = -1.599682593e-08 pk2 = -1.387778781e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.339715233e-01 ldsub = 3.033024110e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.158159998e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.362648555e-9   nfactor = {1.886976015e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.053082948e-7   eta0 = 4.081427101e-01 leta0 = 2.437505465e-8   etab = -1.347621329e-03 letab = 3.799063485e-10   u0 = 7.040683625e-03 lu0 = -5.504378792e-10   ua = -1.613983779e-09 lua = 2.264365708e-16   ub = 2.025147933e-18 lub = -4.321827452e-25   uc = -6.712093967e-11 luc = 1.969220019e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.716932025e+05 lvsat = -1.284569167e-2   a0 = 9.052648244e-01 la0 = -8.651029208e-8   ags = 9.445453886e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.136650759e+00 la2 = -1.014307462e-7   b0 = 1.921756906e-16 lb0 = -5.722511627e-23   b1 = 7.989623218e-20 lb1 = -2.379110054e-26   keta = -4.583734636e-02 lketa = 4.200684472e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.292099820e-01 lpclm = 3.771055897e-07 wpclm = -2.220446049e-22 ppclm = -2.220446049e-28   pdiblc1 = -4.478501477e-01 lpdiblc1 = 2.538472164e-07 wpdiblc1 = -5.551115123e-23 ppdiblc1 = 2.081668171e-28   pdiblc2 = -9.997833428e-03 lpdiblc2 = 5.530975654e-09 wpdiblc2 = -8.673617380e-25 ppdiblc2 = 1.084202172e-31   pdiblcb = 2.653629919e-01 lpdiblcb = -1.647835763e-07 ppdiblcb = 2.775557562e-29   drout = 1.478478000e+00 ldrout = -2.828257447e-7   pscbe1 = 6.876139896e+08 lpscbe1 = 3.345779234e+1   pscbe2 = 2.160022972e-08 lpscbe2 = -3.798272305e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.510363785e+00 lbeta0 = 1.189856830e-7   agidl = 1.490566362e-12 lagidl = -8.164949889e-19   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.471888216e-01 lkt1 = 7.296627166e-9   kt2 = -1.323292858e-02 lkt2 = -1.178601122e-8   at = 3.656378506e+03 lat = 1.912648063e-2   ute = 5.522314189e-01 lute = -4.129603001e-7   ua1 = 5.118987964e-09 lua1 = -1.436452236e-15   ub1 = -4.874445755e-18 lub1 = 1.401068390e-24   uc1 = -2.896530271e-10 luc1 = 5.710342159e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.142 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.290094967e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.382843065e-08 wvth0 = 1.346613551e-07 pvth0 = -4.009878502e-14   k1 = -2.636380082e+00 lk1 = 9.571215026e-07 wk1 = 1.022642203e-06 pk1 = -3.045172819e-13   k2 = 1.690497910e+00 lk2 = -5.131982031e-07 wk2 = -7.325438229e-07 pk2 = 2.181332369e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 7.043277027e+00 ldsub = -1.863680276e-06 wdsub = -3.256127780e-06 pdsub = 9.695934498e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {4.755462865e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.015077562e-07 wvoff = -4.075788729e-07 pvoff = 1.213667989e-13   nfactor = {-1.905268198e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.340614954e-06 wnfactor = 1.513662967e-05 pnfactor = -4.507309900e-12   eta0 = 1.165054841e+01 leta0 = -3.323332303e-06 weta0 = -7.100698036e-06 peta0 = 2.114410358e-12   etab = 1.094859336e+00 letab = -3.260431204e-07 wetab = -6.950155960e-07 petab = 2.069582691e-13   u0 = -9.077133756e-02 lu0 = 2.857553673e-08 wu0 = 6.647842483e-08 pu0 = -1.979561295e-14   ua = -4.960109561e-08 lua = 1.451579880e-14 wua = 3.379667873e-14 pua = -1.006380601e-20   ub = 4.211159248e-17 lub = -1.236892377e-23 wub = -2.884302498e-23 pub = 8.588731764e-30   uc = -5.136100269e-10 luc = 1.526454881e-16 wuc = 3.516977068e-16 puc = -1.047267846e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.624075779e+06 lvsat = 1.415214417e+00 wvsat = 3.142257758e+00 pvsat = -9.356858039e-7   a0 = -1.080760952e+01 la0 = 3.401290866e-06 wa0 = 6.724056742e-06 pa0 = -2.002255996e-12   ags = 2.340909286e+00 lags = -2.484818599e-07 wags = 7.434678650e-15 pags = -2.213859318e-21   a1 = 0.0   a2 = 5.213321537e+00 la2 = -1.315361387e-06 wa2 = -2.712446228e-06 pa2 = 8.076986755e-13   b0 = 0.0   b1 = 0.0   keta = -6.440716365e-01 lketa = 1.823399002e-07 wketa = 3.498951089e-07 pketa = -1.041900161e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.369038781e-01 lpclm = 8.853507505e-11 wpclm = 3.420180887e-08 ppclm = -1.018444364e-14   pdiblc1 = 8.283698114e+00 lpdiblc1 = -2.346189567e-06 wpdiblc1 = -4.910319472e-06 ppdiblc1 = 1.462170381e-12   pdiblc2 = -7.555555349e-02 lpdiblc2 = 2.505242574e-08 wpdiblc2 = 6.872190533e-08 ppdiblc2 = -2.046366536e-14   pdiblcb = -2.880224700e+01 lpdiblcb = 8.490823989e-06 wpdiblcb = 1.990353778e-05 ppdiblcb = -5.926775963e-12   drout = -1.004961910e+00 ldrout = 4.566805746e-07 wdrout = 3.359243500e-12 pdrout = -1.000298735e-18   pscbe1 = 7.998863995e+08 lpscbe1 = 2.587548043e-02 wpscbe1 = 1.004989624e-06 ppscbe1 = -2.992601395e-13   pscbe2 = -7.075382462e-08 lpscbe2 = 2.370245623e-14 wpscbe2 = 5.828269805e-14 ppscbe2 = -1.735513041e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.082166359e+01 lbeta0 = -5.692616161e-07 wbeta0 = -6.523386286e-08 pbeta0 = 1.942501351e-14   agidl = 4.291102656e-08 lagidl = -1.277820358e-14 wagidl = -2.944816462e-14 pagidl = 8.768927220e-21   bgidl = 2.023190686e+09 lbgidl = -2.330572483e+02 wbgidl = 3.730125427e-06 pbgidl = -1.110738754e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -2.394550439e+00 lkt1 = 5.573947328e-07 wkt1 = 1.323447371e-06 pkt1 = -3.940895408e-13   kt2 = 1.813910098e+00 lkt2 = -5.558635261e-07 wkt2 = -1.191865809e-06 pkt2 = 3.549078412e-13   at = -7.173427337e+05 lat = 2.338219913e-01 wat = 6.022892212e-01 pat = -1.793466728e-7   ute = -1.982612902e+01 lute = 5.655205981e-06 wute = 1.135566615e-05 pute = -3.381433489e-12   ua1 = -1.609861027e-08 lua1 = 4.881618078e-15 wua1 = 1.031641450e-14 pua1 = -3.071970328e-21   ub1 = 1.442860349e-17 lub1 = -4.346897099e-24 wub1 = -9.402465310e-24 pub1 = 2.799819108e-30   uc1 = -6.243440599e-10 luc1 = 1.567660439e-16 wuc1 = 1.929610835e-16 puc1 = -5.745898665e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.143 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-07 wmax = 7.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-5.367374994e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.158108050e-07 wvth0 = -3.413306284e-07 pvth0 = 7.341937765e-14   k1 = 4.019487767e+00 lk1 = -6.006337329e-07 wk1 = -1.939749170e-06 pk1 = 3.978744019e-13   k2 = -2.502456178e+00 lk2 = 4.748295569e-07 wk2 = 1.587016031e-06 pk2 = -3.333566399e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -8.951888059e+00 ldsub = 1.912440375e-06 wdsub = 6.176231601e-06 pdsub = -1.266846656e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.387133483e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.393901416e-07 wvoff = 7.733800164e-07 pvoff = -1.586441954e-13   nfactor = {4.510544343e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.890458037e-06 wnfactor = -2.872173896e-05 pnfactor = 5.891718952e-12   eta0 = -1.997826888e+01 leta0 = 4.170574354e-06 weta0 = 1.347356387e-05 peta0 = -2.763845465e-12   etab = -2.004250866e+00 letab = 4.082073326e-07 wetab = 1.318306898e-06 petab = -2.704064022e-13   u0 = 1.833731897e-01 lu0 = -3.639545313e-08 wu0 = -1.183447695e-07 pu0 = 2.396703775e-14   ua = 9.522399237e-08 lua = -1.985037465e-14 wua = -6.412913019e-14 pua = 1.315487114e-20   ub = -8.140158564e-17 lub = 1.694085908e-23 wub = 5.472957941e-23 pub = -1.122673200e-29   uc = 1.000444143e-09 luc = -2.065644166e-16 wuc = -6.671005802e-16 puc = 1.368332766e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.171936802e+07 lvsat = -2.479627430e+00 wvsat = -7.921314468e+00 pvsat = 1.702565125e-6   a0 = 2.025970039e+01 la0 = -3.949354381e-06 wa0 = -1.275888486e-05 pa0 = 2.617242546e-12   ags = 1.250000099e+00 lags = -2.129070609e-14 wags = -1.864231081e-14 pags = 4.003901211e-21   a1 = 0.0   a2 = -7.069993512e+00 la2 = 1.593114983e-06 wa2 = 5.144971027e-06 pa2 = -1.055317997e-12   b0 = 0.0   b1 = 0.0   keta = 9.960422467e-01 lketa = -2.055100268e-07 wketa = -6.639257830e-07 pketa = 1.361917650e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 7.193590291e-01 lpclm = -2.008781671e-08 wpclm = -6.487376155e-08 ppclm = 1.330666259e-14   pdiblc1 = -1.379903529e+01 lpdiblc1 = 2.884003511e-06 wpdiblc1 = 9.313900444e-06 ppdiblc1 = -1.910433880e-12   pdiblc2 = 1.993295169e-01 lpdiblc2 = -4.036277815e-08 wpdiblc2 = -1.303517628e-07 ppdiblc2 = 2.673728493e-14   pdiblcb = 5.623332924e+01 lpdiblcb = -1.169004606e-05 wpdiblcb = -3.775304988e-05 ppdiblcb = 7.743770024e-12   drout = 1.000013454e+00 ldrout = -2.889597866e-12 wdrout = -8.423241937e-12 pdrout = 1.809101786e-18   pscbe1 = 8.000000046e+08 lpscbe1 = -9.837989807e-07 wpscbe1 = -2.519989014e-06 ppscbe1 = 5.412311554e-13   pscbe2 = 1.731557523e-07 lpscbe2 = -3.423147631e-14 wpscbe2 = -1.105506879e-13 ppscbe2 = 2.267576048e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.165899764e+00 lbeta0 = 3.831610131e-08 wbeta0 = 1.237396921e-07 pbeta0 = -2.538120143e-14   agidl = -1.075805654e-07 lagidl = 2.310467391e-14 wagidl = 7.383678152e-14 pagidl = -1.585817609e-20   bgidl = 1.000000369e+09 lbgidl = -7.913546753e-05 wbgidl = -9.353210449e-06 pbgidl = 2.008838654e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 3.228243159e+00 lkt1 = -7.773233828e-07 wkt1 = -2.511240611e-06 pkt1 = 5.151333147e-13   kt2 = -3.486365399e+00 lkt2 = 7.000245032e-07 wkt2 = 2.260731847e-06 pkt2 = -4.637131832e-13   at = 1.754392140e+06 lat = -3.537455950e-01 wat = -1.142422768e+00 pat = 2.343296553e-7   ute = 3.224971247e+01 lute = -6.669581503e-06 wute = -2.153943964e-05 pute = 4.418092552e-12   ua1 = 3.008726929e-08 lua1 = -6.059190749e-15 wua1 = -1.956818090e-14 pua1 = 4.013754832e-21   ub1 = -2.721668834e-17 lub1 = 5.522398298e-24 wub1 = 1.783460617e-23 pub1 = -3.658170405e-30   uc1 = 5.269136021e-10 luc1 = -1.133328078e-16 wuc1 = -3.660087535e-16 puc1 = 7.507440050e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.144 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.145 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124300389e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.583094798e-7   k1 = 4.169979224e-01 lk1 = 2.938540225e-7   k2 = 5.787523347e-02 lk2 = -3.323321159e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 2.964615315e-27   voff = {-1.544415308e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.787950865e-7   nfactor = {1.810230600e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.882834906e-6   eta0 = 0.08   etab = -0.07   u0 = 6.082762501e-03 lu0 = 3.565351435e-8   ua = -6.616112197e-10 lua = -1.158519626e-15   ub = 4.662300295e-20 lub = 1.125904990e-23 pub = 6.162975822e-45   uc = -1.046504257e-10 luc = -2.029966214e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.296000734e+04 lvsat = -2.566918583e-1   a0 = 1.627020626e+00 la0 = -3.268200833e-6   ags = 1.127420605e-01 lags = 1.098496716e-8   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 1.250763844e-07 lb0 = -1.957753127e-12 pb0 = -4.235164736e-34   b1 = -6.804545270e-09 lb1 = 5.623491643e-14   keta = 3.424649349e-02 lketa = -2.182247320e-07 pketa = 2.220446049e-28   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-6   pdiblc1 = 0.39   pdiblc2 = 1.911548633e-03 lpdiblc2 = -1.271810464e-8   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.857143290e-09 lpscbe2 = 2.412713055e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.810749375e+01 lbeta0 = -3.630149605e-4   agidl = 2.814705940e-09 lagidl = -1.833265859e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.444100755e-01 lkt1 = 1.234958073e-7   kt2 = -6.524363936e-02 lkt2 = 1.342727668e-7   at = 7.717891133e+04 lat = -1.240739019e-1   ute = 5.643158221e-01 lute = -1.297684100e-05 wute = 1.110223025e-22 pute = 4.440892099e-27   ua1 = 3.780637815e-09 lua1 = -3.388951696e-14 pua1 = -2.646977960e-35   ub1 = -2.653212355e-18 lub1 = 2.855429361e-23 pub1 = 1.232595164e-44   uc1 = -9.464587252e-11 luc1 = 1.300235988e-15 puc1 = 8.271806126e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.146 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140859468e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.504573657e-8   k1 = 4.604519148e-01 lk1 = -5.585393079e-8   k2 = 1.358353148e-02 lk2 = 2.411753606e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.414495418e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.214258093e-7   nfactor = {9.948645590e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.679047535e-6   eta0 = 0.08   etab = -0.07   u0 = 9.506801114e-03 lu0 = 8.097621998e-9   ua = -9.746330556e-10 lua = 1.360609680e-15   ub = 1.472299687e-18 lub = -2.144752731e-25   uc = -1.070061023e-10 luc = -1.341706802e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.345534345e+04 lvsat = -1.924496188e-2   a0 = 1.168891106e+00 la0 = 4.187224649e-7   ags = 4.434987157e-02 lags = 5.613899157e-7   a1 = 0.0   a2 = 0.8   b0 = -8.806443456e-08 lb0 = -2.424437724e-13   b1 = 3.575823691e-09 lb1 = -2.730395738e-14 wb1 = -1.240770919e-30 pb1 = 4.963083675e-36   keta = 7.542872474e-03 lketa = -3.319998307e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -4.142606150e-01 lpclm = 4.468282376e-06 ppclm = 1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 2.312663529e-04 lpdiblc2 = 8.044290883e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.465165627e-08 lpscbe2 = -2.250580619e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.011943750e-10 lalpha0 = -8.143895613e-16   alpha1 = 2.011943750e-10 lalpha1 = -8.143895613e-16   beta0 = -2.432248125e+01 lbeta0 = 2.198851815e-04 pbeta0 = -1.136868377e-25   agidl = 6.955865393e-10 lagidl = -1.278462449e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.136981111e-01 lkt1 = -1.236671723e-7   kt2 = -3.845308193e-02 lkt2 = -8.133161144e-8   at = 2.206495351e+04 lat = 3.194708301e-1   ute = -1.923673091e+00 lute = 7.045933977e-6   ua1 = -2.981113444e-09 lua1 = 2.052753578e-14 wua1 = 8.271806126e-31 pua1 = 3.308722450e-36   ub1 = 2.942842689e-18 lub1 = -1.648149826e-23 wub1 = 1.540743956e-39 pub1 = 6.162975822e-45   uc1 = 5.577709848e-10 luc1 = -3.950268087e-15 wuc1 = 1.033975766e-31 puc1 = 4.135903063e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.147 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.145429258e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.548256636e-9   k1 = 3.846063128e-01 lk1 = 2.511520008e-7   k2 = 4.228702503e-02 lk2 = -9.206774752e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.671662398e-01 ldsub = -1.243339826e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.160605222e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.865677060e-8   nfactor = {2.216222452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.647344113e-7   eta0 = 1.613990562e-01 leta0 = -3.294850649e-7   etab = -1.411601813e-01 letab = 2.880404027e-7   u0 = 1.273220293e-02 lu0 = -4.958078823e-9   ua = -3.083681764e-10 lua = -1.336280642e-15   ub = 1.131103764e-18 lub = 1.166609054e-24   uc = -1.341261632e-10 luc = 1.084341980e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.419147855e+04 lvsat = -1.031801711e-1   a0 = 1.402304588e+00 la0 = -5.260827937e-7   ags = -4.704625846e-02 lags = 9.313408859e-7   a1 = 0.0   a2 = 0.8   b0 = -1.959803237e-07 lb0 = 1.943754660e-13 wb0 = 2.117582368e-28   b1 = -3.047654999e-09 lb1 = -4.936059274e-16   keta = 2.300377997e-02 lketa = -6.590227314e-08 wketa = -1.387778781e-23   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.049877559e-01 lpclm = 3.425943017e-7   pdiblc1 = 0.39   pdiblc2 = 4.184058358e-04 lpdiblc2 = 4.693056786e-11   pdiblcb = -4.297775000e-01 lpdiblcb = 8.288932451e-7   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.707934004e-09 lpscbe2 = 1.553044224e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.023887500e-10 lalpha0 = 4.144466225e-16   alpha1 = -1.023887500e-10 lalpha1 = 4.144466225e-16   beta0 = 5.501572660e+01 lbeta0 = -1.012580327e-4   agidl = -7.892498222e-11 lagidl = 1.856585925e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.354240898e-01 lkt1 = -3.572529886e-8   kt2 = -6.326714526e-02 lkt2 = 1.911013376e-8   at = 1.633938954e+05 lat = -2.525969275e-1   ute = -9.045128663e-02 lute = -3.745354128e-7   ua1 = 2.896511406e-09 lua1 = -3.263767152e-15   ub1 = -1.914119324e-18 lub1 = 3.178391148e-24   uc1 = -8.826429466e-10 luc1 = 1.880203415e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.148 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.156253754e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.561787663e-8   k1 = 5.064465886e-01 lk1 = 1.650529987e-9   k2 = -2.574283335e-03 lk2 = -2.018817928e-10   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.600000205e-01 ldsub = -2.145607514e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.095058695e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.234316656e-9   nfactor = {2.507545012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.612974670e-7   eta0 = -5.123858625e-01 leta0 = 1.050274847e-06 weta0 = -9.454242944e-23 peta0 = -3.868433351e-28   etab = 2.826599494e-04 letab = -1.602711478e-9   u0 = 1.299327309e-02 lu0 = -5.492691778e-9   ua = -3.839322797e-10 lua = -1.181542360e-15   ub = 1.453484210e-18 lub = 5.064464363e-25   uc = -1.205586833e-10 luc = 8.065105179e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.493717597e+04 lvsat = 3.863705835e-2   a0 = 1.028226064e+00 la0 = 2.399458559e-7   ags = 2.437725462e-01 lags = 3.358094083e-7   a1 = 0.0   a2 = 0.8   b0 = -6.697383500e-09 lb0 = -1.932334070e-13   b1 = -6.829548739e-09 lb1 = 7.250861527e-15   keta = -1.770930147e-02 lketa = 1.746895719e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.234158669e-01 lpclm = -3.094748232e-7   pdiblc1 = 3.959313076e-01 lpdiblc1 = -1.214598339e-8   pdiblc2 = 4.531883283e-04 lpdiblc2 = -2.429615072e-11   pdiblcb = 1.845550000e-01 lpdiblcb = -4.291214901e-07 wpdiblcb = 5.551115123e-23 ppdiblcb = -2.220446049e-28   drout = 3.752086697e-01 ldrout = 3.784110665e-7   pscbe1 = 800000000.0   pscbe2 = 9.776711087e-09 lpscbe2 = -6.355707662e-16 wpscbe2 = 1.323488980e-29   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.621328974e+00 lbeta0 = 1.938354859e-6   agidl = 4.019000103e-10 lagidl = 8.719645261e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.254238063e-01 lkt1 = -5.620362931e-8   kt2 = -5.956764875e-02 lkt2 = 1.153439730e-8   at = 2.776234628e+04 lat = 2.514596790e-2   ute = 5.384763382e-01 lute = -1.662437680e-06 pute = -4.440892099e-28   ua1 = 3.118603033e-09 lua1 = -3.718560834e-15   ub1 = -1.637022257e-18 lub1 = 2.610958703e-24   uc1 = 2.633427840e-12 luc1 = 6.735658696e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.149 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.394755713e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.655142663e-07 wvth0 = 1.180478678e-07 pvth0 = -1.236876047e-13   k1 = -2.808768743e-01 lk1 = 8.265883714e-07 wk1 = 5.007202577e-07 pk1 = -5.246421680e-13   k2 = 4.766831099e-01 lk2 = -5.023557970e-07 wk2 = -3.010962502e-07 pk2 = 3.154811236e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 7.352065134e+00 ldsub = -7.430888546e-06 wdsub = -4.553830192e-06 pdsub = 4.771389430e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {2.743186355e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.017049041e-07 wvoff = -3.023171542e-07 pvoff = 3.167603562e-13   nfactor = {-9.396071851e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.161101469e-05 wnfactor = 6.776042395e-06 pnfactor = -7.099767821e-12   eta0 = -4.145574603e+00 leta0 = 4.857039180e-06 weta0 = 2.975341014e-06 peta0 = -3.117487931e-12   etab = -5.536146206e-03 letab = 4.494088141e-09 wetab = 2.315645993e-09 petab = -2.426275980e-15   u0 = 1.695738889e-02 lu0 = -9.646193205e-09 wu0 = -4.661839959e-09 pu0 = 4.884559363e-15   ua = 5.693188735e-09 lua = -7.548997831e-15 wua = -4.800685983e-15 pua = 5.030038756e-21   ub = -9.207515841e-18 lub = 1.167677577e-23 wub = 7.578777911e-24 pub = -7.940854026e-30   uc = -2.377444434e-10 luc = 2.034353615e-16 wuc = 1.148778865e-16 puc = -1.203661776e-22   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -5.273346598e+05 lvsat = 6.068159311e-01 wvsat = 3.012579331e-01 pvsat = -3.156505308e-7   a0 = 5.676882140e+00 la0 = -4.630799763e-06 wa0 = -2.456513125e-06 pa0 = 2.573873039e-12   ags = -1.869811236e-01 lags = 7.871423346e-07 wags = -3.954223615e-16 pags = 4.143139165e-22   a1 = 0.0   a2 = -4.198763207e+00 la2 = 5.237579119e-06 wa2 = 3.074786438e-06 pa2 = -3.221684360e-12   b0 = -4.005015170e-07 lb0 = 2.193847190e-13 wb0 = 5.871242755e-22 pb0 = -6.151741951e-28   b1 = 1.900621935e-10 lb1 = -1.041113178e-16 wb1 = 2.440943813e-25 pb1 = -2.557560770e-31   keta = -1.677644320e-02 lketa = 1.649153163e-08 wketa = 3.589580655e-08 pketa = -3.761072871e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.178756718e+00 lpclm = -4.768114584e-06 wpclm = -2.498815450e-06 ppclm = 2.618196358e-12   pdiblc1 = 1.359745187e+00 lpdiblc1 = -1.022006071e-06 wpdiblc1 = -3.635401056e-07 ppdiblc1 = 3.809082342e-13   pdiblc2 = 8.202531298e-03 lpdiblc2 = -8.143863980e-09 wpdiblc2 = -4.714650707e-09 ppdiblc2 = 4.939893145e-15   pdiblcb = -2.426893159e+00 lpdiblcb = 2.307088604e-06 wpdiblcb = 1.268801299e-06 ppdiblcb = -1.329418281e-12   drout = -4.247639314e+00 ldrout = 5.222115612e-06 wdrout = 3.013598690e-06 pdrout = -3.157573367e-12   pscbe1 = -5.566216108e+09 lpscbe1 = 6.670362082e+03 wpscbe1 = 4.086152313e+03 ppscbe1 = -4.281368240e-3   pscbe2 = 6.713559027e-07 lpscbe2 = -6.938217082e-13 wpscbe2 = -4.251347042e-13 ppscbe2 = 4.454455147e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.959682000e-01 lbeta0 = 5.736917244e-06 wbeta0 = 1.910901841e-06 pbeta0 = -2.002195176e-12   agidl = 1.219645083e-08 lagidl = -1.148607096e-14 wagidl = -6.114393250e-15 pagidl = 6.406508388e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 1.069284623e-01 lkt1 = -6.139890275e-07 wkt1 = -3.346282048e-07 pkt1 = 3.506150673e-13   kt2 = -3.245689587e-01 lkt2 = 2.891961448e-07 wkt2 = 1.659802832e-07 pkt2 = -1.739099913e-13   at = 5.020849190e+05 lat = -4.718373658e-01 wat = -2.773171810e-01 pat = 2.905660093e-7   ute = -2.364262007e+00 lute = 1.378978990e-06 wute = 2.473124173e-07 pute = -2.591277680e-13   ua1 = -1.238102154e-08 lua1 = 1.252155831e-14 wua1 = 5.563139867e-15 pua1 = -5.828918874e-21   ub1 = 1.958846686e-17 lub1 = -1.962857816e-23 wub1 = -9.708231753e-24 pub1 = 1.017204253e-29   uc1 = 1.585502296e-09 luc1 = -1.591133842e-15 wuc1 = -7.902943775e-16 puc1 = 8.280506914e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.150 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-7.126737840e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.081131622e-07 wvth0 = -2.360957356e-07 pvth0 = 7.030340768e-14   k1 = 2.002630472e+00 lk1 = -4.242598650e-07 wk1 = -1.001440515e-06 pk1 = 2.982039495e-13   k2 = -9.257220738e-01 lk2 = 2.658467025e-07 wk2 = 6.021925004e-07 pk2 = -1.793178718e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -1.454897043e+01 ldsub = 4.565951210e-06 wdsub = 9.107660384e-06 pdsub = -2.712033571e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.166152211e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.873490138e-07 wvoff = 6.046343083e-07 pvoff = -1.800449812e-13   nfactor = {2.318751543e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.237459828e-06 wnfactor = -1.355208479e-05 pnfactor = 4.035472049e-12   eta0 = 9.761149206e+00 leta0 = -2.760716455e-06 weta0 = -5.950682029e-06 peta0 = 1.771964341e-12   etab = 5.931628985e-03 letab = -1.787672414e-09 wetab = -4.631291985e-09 petab = 1.379082971e-15   u0 = -7.613844783e-03 lu0 = 3.813314318e-09 wu0 = 9.323679919e-09 pu0 = -2.776358788e-15   ua = -1.670497569e-08 lua = 4.720156687e-15 wua = 9.601371966e-15 pua = -2.859048537e-21   ub = 2.584909238e-17 lub = -7.526357802e-24 wub = -1.515755582e-23 pub = 4.513541185e-30   uc = 2.939985467e-10 luc = -8.784015487e-17 wuc = -2.297557731e-16 puc = 6.841552532e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.118699744e+06 lvsat = -2.948405647e-01 wvsat = -6.025158662e-01 pvsat = 1.794141621e-7   a0 = -6.816802361e+00 la0 = 2.212928264e-06 wa0 = 4.913026249e-06 pa0 = -1.462976391e-12   ags = 9.445453874e-01 lags = 1.673204001e-07 wags = 7.908482758e-16 pags = -2.354934026e-22   a1 = 0.0   a2 = 1.080226468e+01 la2 = -2.979608931e-06 wa2 = -6.149572875e-06 pa2 = 1.831189063e-12   b0 = 2.037805400e-15 lb0 = -6.068075029e-22 wb0 = -1.174248681e-21 pb0 = 3.496619010e-28   b1 = 8.472089932e-19 lb1 = -2.522776580e-25 wb1 = -4.881889326e-25 pb1 = 1.453704594e-31   keta = 6.700138717e-02 lketa = -2.939986940e-08 wketa = -7.179161311e-08 pketa = 2.137774759e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -8.484254839e+00 lpclm = 2.716141572e-06 wpclm = 4.997630900e-06 ppclm = -1.488169541e-12   pdiblc1 = -1.590641160e+00 lpdiblc1 = 5.941418100e-07 wpdiblc1 = 7.270802113e-07 ppdiblc1 = -2.165063099e-13   pdiblc2 = -2.481837281e-02 lpdiblc2 = 9.944161769e-09 wpdiblc2 = 9.429301414e-09 ppdiblc2 = -2.807810229e-15   pdiblcb = 4.253849263e+00 lpdiblcb = -1.352455076e-06 wpdiblcb = -2.537602597e-06 ppdiblcb = 7.556346134e-13   drout = 1.095174778e+01 ldrout = -3.103728654e-06 wdrout = -6.027197380e-06 pdrout = 1.794748700e-12   pscbe1 = 1.353246402e+10 lpscbe1 = -3.791417426e+03 wpscbe1 = -8.172304626e+03 ppscbe1 = 2.433508010e-3   pscbe2 = -1.314813859e-06 lpscbe2 = 3.941524329e-13 wpscbe2 = 8.502694085e-13 ppscbe2 = -2.531889731e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.451729786e+01 lbeta0 = -1.669729112e-06 wbeta0 = -3.821803682e-06 pbeta0 = 1.138037591e-12   agidl = -1.921914986e-08 lagidl = 5.722609708e-15 wagidl = 1.222878650e-14 pagidl = -3.641426900e-21   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.599095060e+00 lkt1 = 3.205280072e-07 wkt1 = 6.692564096e-07 pkt1 = -1.992878274e-13   kt2 = 5.085273200e-01 lkt2 = -1.671531692e-07 wkt2 = -3.319605665e-07 pkt2 = 9.884955768e-14   at = -8.680922319e+05 lat = 2.787114231e-01 wat = 5.546343619e-01 pat = -1.651562471e-7   ute = 1.329659833e+00 lute = -6.444590460e-07 wute = -4.946248345e-07 pute = 1.472869101e-13   ua1 = 2.260675930e-08 lua1 = -6.643873346e-15 wua1 = -1.112627973e-14 pua1 = 3.313127948e-21   ub1 = -3.539234411e-17 lub1 = 1.048853557e-23 wub1 = 1.941646351e-23 pub1 = -5.781737421e-30   uc1 = -2.773949251e-09 luc1 = 7.968647296e-16 wuc1 = 1.580588755e-15 puc1 = -4.706598165e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.151 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.078440484e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.030169421e-10   k1 = -1.029038416e+00 lk1 = 4.784953380e-7   k2 = 5.391194458e-01 lk2 = -1.703464810e-07 wk2 = -1.110223025e-22 pk2 = 8.326672685e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.925446141e+00 ldsub = -3.397181839e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.650673151e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.074904104e-8   nfactor = {4.738371709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.437660579e-7   eta0 = 4.900000008e-01 leta0 = -8.645884009e-17   etab = 2.466001640e-03 letab = -7.556952310e-10 wetab = -2.168404345e-25 petab = 5.421010862e-32   u0 = 1.371637263e-02 lu0 = -2.538291171e-9   ua = 3.518959235e-09 lua = -1.302025535e-15 pua = -8.271806126e-37   ub = -3.222538750e-18 lub = 1.130447157e-24   uc = 3.917214497e-11 luc = -1.195922309e-17 wuc = -2.261821987e-32 puc = -4.038967835e-39   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.147794778e+05 lvsat = -5.545320730e-2   a0 = -2.390484591e-01 la0 = 2.542375959e-7   ags = 2.340909298e+00 lags = -2.484818634e-7   a1 = 0.0   a2 = 9.500241430e-01 la2 = -4.585800563e-8   b0 = 0.0   b1 = 0.0   keta = -9.412270452e-02 lketa = 1.857885700e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.906606977e-01 lpclm = -1.591890189e-8   pdiblc1 = 5.658853163e-01 lpdiblc1 = -4.801786142e-8   pdiblc2 = 3.245835548e-02 lpdiblc2 = -7.111415999e-9   pdiblcb = 2.481212150e+00 lpdiblcb = -8.246080592e-07 ppdiblcb = -4.440892099e-28   drout = -1.004956630e+00 ldrout = 4.566790024e-7   pscbe1 = 7.998864011e+08 lpscbe1 = 2.587501007e-2   pscbe2 = 2.085222168e-08 lpscbe2 = -3.575534212e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.071913202e+01 lbeta0 = -5.387302792e-7   agidl = -3.374235138e-09 lagidl = 1.004390227e-15 wagidl = 7.431700816e-31 pagidl = -2.310289601e-37   bgidl = 2.023190692e+09 lbgidl = -2.330572500e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.144171377e-01 lkt1 = -6.201696101e-8   kt2 = -5.940939655e-02 lkt2 = 1.964186534e-9   at = 2.293075782e+05 lat = -4.806680536e-02 pat = 5.820766091e-23   ute = -1.977818730e+00 lute = 3.404253830e-7   ua1 = 1.162523927e-10 lua1 = 5.323734908e-17   ub1 = -3.497561515e-19 lub1 = 5.372894288e-26   uc1 = -3.210567629e-10 luc1 = 6.645466902e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.152 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 7.0e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.056996260e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.386059844e-09 wvth0 = -1.032535659e-08 pvth0 = 2.527389159e-15   k1 = 5.145077898e-04 lk1 = 2.621990477e-07 wk1 = 6.172502245e-07 pk1 = -1.510874237e-13   k2 = 1.919386185e+00 lk2 = -5.209150912e-07 wk2 = -1.226301579e-06 pk2 = 3.001679690e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 3.844660440e+00 ldsub = -8.348487499e-07 wdsub = -1.965342043e-06 pdsub = 4.810665986e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {2.191938413e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.056088209e-07 wvoff = -2.486168299e-07 pvoff = 6.085518453e-14   nfactor = {-1.455019015e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.922080650e-06 wnfactor = 9.233084105e-06 pnfactor = -2.260028162e-12   eta0 = 8.006603801e+00 leta0 = -1.839876695e-06 weta0 = -4.331307640e-06 peta0 = 1.060195827e-12   etab = 7.271532304e-01 letab = -1.781974130e-07 wetab = -4.194997933e-07 petab = 1.026830619e-13   u0 = -5.265406258e-02 lu0 = 1.351808660e-08 wu0 = 3.182332126e-08 pu0 = -7.789553461e-15   ua = -3.797354532e-08 lua = 8.757125518e-15 wua = 2.061540561e-14 pua = -5.046135908e-21   ub = 3.227294475e-17 lub = -7.473588830e-24 wub = -1.759379441e-23 pub = 4.306521026e-30   uc = -3.817241980e-10 luc = 9.017310196e-17 wuc = 2.122791475e-16 puc = -5.196062833e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -8.436272656e+06 lvsat = 2.082446825e+00 wvsat = 4.902349107e+00 pvsat = -1.199972503e-6   a0 = -6.240775311e+00 la0 = 1.742285323e-06 wa0 = 4.101565791e-06 pa0 = -1.003960767e-12   ags = 1.250000069e+00 lags = -1.481563316e-14 wags = 4.728804015e-16 pags = -1.157474117e-22   a1 = 0.0   a2 = 3.589892035e+00 la2 = -6.954542838e-07 wa2 = -1.637189274e-06 pa2 = 4.007430046e-13   b0 = 0.0   b1 = 0.0   keta = -3.829446891e-01 lketa = 9.066189232e-08 wketa = 2.134298332e-07 pketa = -5.224228742e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 5.849462766e-01 lpclm = 8.769237392e-09 wpclm = 2.064393284e-08 ppclm = -5.053118660e-15   pdiblc1 = 5.498469336e+00 lpdiblc1 = -1.258974931e-06 wpdiblc1 = -2.963789519e-06 ppdiblc1 = 7.254615795e-13   pdiblc2 = -7.074685827e-02 lpdiblc2 = 1.761987926e-08 wpdiblc2 = 4.147946957e-08 ppdiblc2 = -1.015313716e-14   pdiblcb = -2.198736783e+01 lpdiblcb = 5.103143937e-06 wpdiblcb = 1.201346066e-05 ppdiblcb = -2.940594833e-12   drout = 1.000000244e+00 ldrout = -5.338899456e-14 wdrout = -1.885381806e-14 pdrout = 4.614943094e-21   pscbe1 = 8.000000019e+08 lpscbe1 = -4.523258209e-07 wpscbe1 = -8.297042847e-07 ppscbe1 = 2.030906677e-13   pscbe2 = -5.589464667e-08 lpscbe2 = 1.494332029e-14 wpscbe2 = 3.517850560e-14 ppscbe2 = -8.610818709e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.422268254e+00 lbeta0 = -1.672361504e-08 wbeta0 = -3.937014558e-08 pbeta0 = 9.636827385e-15   agidl = 7.989983812e-08 lagidl = -1.930405833e-14 wagidl = -4.544425060e-14 pagidl = 1.112361644e-20   bgidl = 1.000000335e+09 lbgidl = -7.134772491e-05 wbgidl = 1.203543854e-05 pbgidl = -2.945976257e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -1.987654248e+00 lkt1 = 3.429210134e-07 wkt1 = 8.072802284e-07 pkt1 = -1.976020179e-13   kt2 = 1.197654862e+00 lkt2 = -3.055871201e-07 wkt2 = -7.193917319e-07 pkt2 = 1.760891112e-13   at = -6.125982525e+05 lat = 1.544232256e-01 wat = 3.635322633e-01 pat = -8.898360975e-8   ute = -1.237793774e+01 lute = 2.911522181e-06 wute = 6.854099510e-06 pute = -1.677712208e-12   ua1 = -1.045613264e-08 lua1 = 2.645066267e-15 wua1 = 6.226828791e-15 pua1 = -1.524172017e-21   ub1 = 9.734902815e-18 lub1 = -2.410733393e-24 wub1 = -5.675178578e-24 pub1 = 1.389141836e-30   uc1 = -2.314214543e-10 luc1 = 4.947403433e-17 wuc1 = 1.164682761e-16 puc1 = -2.850852229e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.153 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.154 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124300389e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.583094798e-7   k1 = 4.169979224e-01 lk1 = 2.938540225e-7   k2 = 5.787523347e-02 lk2 = -3.323321159e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 6.776263578e-27 pcit = 1.897353802e-31   voff = {-1.544415308e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.787950865e-7   nfactor = {1.810230600e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.882834906e-6   eta0 = 0.08   etab = -0.07   u0 = 6.082762501e-03 lu0 = 3.565351435e-8   ua = -6.616112197e-10 lua = -1.158519626e-15   ub = 4.662300295e-20 lub = 1.125904990e-23   uc = -1.046504257e-10 luc = -2.029966214e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.296000734e+04 lvsat = -2.566918583e-1   a0 = 1.627020626e+00 la0 = -3.268200833e-6   ags = 1.127420605e-01 lags = 1.098496716e-8   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 1.250763844e-07 lb0 = -1.957753127e-12 wb0 = 2.117582368e-28 pb0 = -5.082197684e-33   b1 = -6.804545270e-09 lb1 = 5.623491643e-14   keta = 3.424649349e-02 lketa = -2.182247320e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 wpclm = -1.110223025e-22 ppclm = -1.776356839e-27   pdiblc1 = 0.39   pdiblc2 = 1.911548633e-03 lpdiblc2 = -1.271810464e-8   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.857143290e-09 lpscbe2 = 2.412713055e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.810749375e+01 lbeta0 = -3.630149605e-4   agidl = 2.814705940e-09 lagidl = -1.833265859e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.444100755e-01 lkt1 = 1.234958073e-7   kt2 = -6.524363936e-02 lkt2 = 1.342727668e-7   at = 7.717891133e+04 lat = -1.240739019e-01 wat = 4.656612873e-16   ute = 5.643158221e-01 lute = -1.297684100e-05 wute = 8.881784197e-22 pute = -2.131628207e-26   ua1 = 3.780637815e-09 lua1 = -3.388951696e-14 pua1 = -1.058791184e-34   ub1 = -2.653212355e-18 lub1 = 2.855429361e-23 wub1 = 1.232595164e-38   uc1 = -9.464587252e-11 luc1 = 1.300235988e-15 puc1 = -1.654361225e-36   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.155 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140859468e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.504573657e-8   k1 = 4.604519148e-01 lk1 = -5.585393079e-8   k2 = 1.358353148e-02 lk2 = 2.411753606e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.414495418e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.214258093e-7   nfactor = {9.948645590e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.679047535e-6   eta0 = 0.08   etab = -0.07   u0 = 9.506801114e-03 lu0 = 8.097621998e-9   ua = -9.746330556e-10 lua = 1.360609680e-15   ub = 1.472299687e-18 lub = -2.144752731e-25   uc = -1.070061023e-10 luc = -1.341706802e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.345534345e+04 lvsat = -1.924496188e-2   a0 = 1.168891106e+00 la0 = 4.187224649e-7   ags = 4.434987157e-02 lags = 5.613899157e-7   a1 = 0.0   a2 = 0.8   b0 = -8.806443456e-08 lb0 = -2.424437724e-13   b1 = 3.575823691e-09 lb1 = -2.730395738e-14 wb1 = 4.963083675e-30 pb1 = -2.646977960e-35   keta = 7.542872474e-03 lketa = -3.319998307e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -4.142606150e-01 lpclm = 4.468282376e-06 ppclm = 1.421085472e-26   pdiblc1 = 0.39   pdiblc2 = 2.312663529e-04 lpdiblc2 = 8.044290883e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.465165627e-08 lpscbe2 = -2.250580619e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.011943750e-10 lalpha0 = -8.143895613e-16   alpha1 = 2.011943750e-10 lalpha1 = -8.143895613e-16   beta0 = -2.432248125e+01 lbeta0 = 2.198851815e-04 wbeta0 = 5.684341886e-20 pbeta0 = 4.547473509e-25   agidl = 6.955865393e-10 lagidl = -1.278462449e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.136981111e-01 lkt1 = -1.236671723e-7   kt2 = -3.845308193e-02 lkt2 = -8.133161144e-8   at = 2.206495351e+04 lat = 3.194708301e-1   ute = -1.923673091e+00 lute = 7.045933977e-6   ua1 = -2.981113444e-09 lua1 = 2.052753578e-14 wua1 = -3.308722450e-30 pua1 = 3.970466940e-35   ub1 = 2.942842689e-18 lub1 = -1.648149826e-23 pub1 = -4.930380658e-44   uc1 = 5.577709848e-10 luc1 = -3.950268087e-15 wuc1 = 8.271806126e-31 puc1 = -9.926167351e-36   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.156 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.145429258e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.548256636e-9   k1 = 3.846063128e-01 lk1 = 2.511520008e-7   k2 = 4.228702503e-02 lk2 = -9.206774752e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.671662398e-01 ldsub = -1.243339826e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.160605222e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.865677060e-8   nfactor = {2.216222452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.647344113e-7   eta0 = 1.613990562e-01 leta0 = -3.294850649e-7   etab = -1.411601813e-01 letab = 2.880404027e-7   u0 = 1.273220293e-02 lu0 = -4.958078823e-9   ua = -3.083681764e-10 lua = -1.336280642e-15   ub = 1.131103764e-18 lub = 1.166609054e-24   uc = -1.341261632e-10 luc = 1.084341980e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.419147855e+04 lvsat = -1.031801711e-1   a0 = 1.402304588e+00 la0 = -5.260827937e-7   ags = -4.704625846e-02 lags = 9.313408859e-7   a1 = 0.0   a2 = 0.8   b0 = -1.959803238e-07 lb0 = 1.943754660e-13   b1 = -3.047654999e-09 lb1 = -4.936059274e-16   keta = 2.300377997e-02 lketa = -6.590227314e-08 wketa = -5.551115123e-23 pketa = -1.110223025e-28   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.049877559e-01 lpclm = 3.425943017e-7   pdiblc1 = 0.39   pdiblc2 = 4.184058358e-04 lpdiblc2 = 4.693056786e-11   pdiblcb = -4.297775000e-01 lpdiblcb = 8.288932451e-7   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.707934004e-09 lpscbe2 = 1.553044224e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.023887500e-10 lalpha0 = 4.144466225e-16   alpha1 = -1.023887500e-10 lalpha1 = 4.144466225e-16   beta0 = 5.501572660e+01 lbeta0 = -1.012580327e-4   agidl = -7.892498222e-11 lagidl = 1.856585925e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.354240898e-01 lkt1 = -3.572529886e-8   kt2 = -6.326714526e-02 lkt2 = 1.911013376e-8   at = 1.633938953e+05 lat = -2.525969275e-1   ute = -9.045128663e-02 lute = -3.745354128e-7   ua1 = 2.896511406e-09 lua1 = -3.263767152e-15   ub1 = -1.914119324e-18 lub1 = 3.178391148e-24   uc1 = -8.826429466e-10 luc1 = 1.880203415e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.157 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.156253754e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.561787663e-8   k1 = 5.064465886e-01 lk1 = 1.650529987e-9   k2 = -2.574283335e-03 lk2 = -2.018817928e-10   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.600000205e-01 ldsub = -2.145607425e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.095058695e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.234316656e-9   nfactor = {2.507545012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.612974670e-7   eta0 = -5.123858625e-01 leta0 = 1.050274847e-06 weta0 = 8.881784197e-22 peta0 = -1.665334537e-27   etab = 2.826599494e-04 letab = -1.602711478e-9   u0 = 1.299327309e-02 lu0 = -5.492691778e-9   ua = -3.839322797e-10 lua = -1.181542360e-15   ub = 1.453484210e-18 lub = 5.064464363e-25   uc = -1.205586833e-10 luc = 8.065105179e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.493717597e+04 lvsat = 3.863705835e-2   a0 = 1.028226064e+00 la0 = 2.399458559e-7   ags = 2.437725462e-01 lags = 3.358094083e-7   a1 = 0.0   a2 = 0.8   b0 = -6.697383500e-09 lb0 = -1.932334070e-13   b1 = -6.829548739e-09 lb1 = 7.250861527e-15   keta = -1.770930147e-02 lketa = 1.746895719e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.234158669e-01 lpclm = -3.094748232e-7   pdiblc1 = 3.959313076e-01 lpdiblc1 = -1.214598339e-8   pdiblc2 = 4.531883283e-04 lpdiblc2 = -2.429615072e-11   pdiblcb = 1.845550000e-01 lpdiblcb = -4.291214901e-07 ppdiblcb = -4.440892099e-28   drout = 3.752086697e-01 ldrout = 3.784110665e-7   pscbe1 = 800000000.0   pscbe2 = 9.776711087e-09 lpscbe2 = -6.355707662e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.621328974e+00 lbeta0 = 1.938354859e-6   agidl = 4.019000103e-10 lagidl = 8.719645261e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.254238063e-01 lkt1 = -5.620362931e-8   kt2 = -5.956764875e-02 lkt2 = 1.153439730e-8   at = 2.776234628e+04 lat = 2.514596790e-2   ute = 5.384763382e-01 lute = -1.662437680e-06 pute = 3.552713679e-27   ua1 = 3.118603033e-09 lua1 = -3.718560834e-15   ub1 = -1.637022257e-18 lub1 = 2.610958703e-24 wub1 = -3.081487911e-39 pub1 = -3.081487911e-45   uc1 = 2.633427840e-12 luc1 = 6.735658696e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.158 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.189894012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.086529730e-8   k1 = 5.880791324e-01 lk1 = -8.388200862e-8   k2 = -4.584297371e-02 lk2 = 4.513397027e-08 wk2 = -8.326672685e-23 pk2 = 5.551115123e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.507070000e-01 ldsub = 8.494385269e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.503262196e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.800485898e-8   nfactor = {2.363154285e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.100084730e-07 wnfactor = -1.421085472e-20   eta0 = 1.017868271e+00 leta0 = -5.530871778e-7   etab = -1.517546071e-03 letab = 2.834993852e-10   u0 = 8.867175292e-03 lu0 = -1.169469657e-9   ua = -2.637979932e-09 lua = 1.180192418e-15   ub = 3.944787243e-18 lub = -2.103878599e-24   uc = -3.838396610e-11 luc = -5.449562538e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.527989752e+03 lvsat = 5.903217237e-2   a0 = 1.413819476e+00 la0 = -1.640692811e-7   ags = -1.869811243e-01 lags = 7.871423354e-7   a1 = 0.0   a2 = 1.137258461e+00 la2 = -3.533709843e-07 wa2 = -7.105427358e-21   b0 = -4.005015160e-07 lb0 = 2.193847179e-13   b1 = 1.900621939e-10 lb1 = -1.041113183e-16   keta = 4.551757475e-02 lketa = -4.877858303e-08 wketa = 6.938893904e-23 pketa = 8.326672685e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 8.422820869e-01 lpclm = -2.244648769e-7   pdiblc1 = 7.288532800e-01 lpdiblc1 = -3.609733030e-7   pdiblc2 = 2.066929197e-05 lpdiblc2 = 4.288864826e-10   pdiblcb = -0.225   drout = 9.821963946e-01 ldrout = -2.575754971e-07 wdrout = -7.105427358e-21   pscbe1 = 1.524942164e+09 lpscbe1 = -7.595762759e+2   pscbe2 = -6.642801811e-08 lpscbe2 = 7.920983936e-14 wpscbe2 = -2.117582368e-28 ppscbe2 = 5.293955920e-35   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.312170425e+00 lbeta0 = 2.262283457e-6   agidl = 1.585458645e-09 lagidl = -3.681386223e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.737893819e-01 lkt1 = -5.527388326e-9   kt2 = -3.652476254e-02 lkt2 = -1.260936280e-8   at = 2.082532054e+04 lat = 3.241441004e-2   ute = -1.935073039e+00 lute = 9.292855189e-7   ua1 = -2.726681161e-09 lua1 = 2.405981813e-15 wua1 = 3.308722450e-30 pua1 = 3.308722450e-36   ub1 = 2.740683756e-18 lub1 = -1.975892216e-24 pub1 = 6.162975822e-45   uc1 = 2.140158506e-10 luc1 = -1.541246310e-16 puc1 = 4.135903063e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.159 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.122397186e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.389222392e-8   k1 = 2.647184581e-01 lk1 = 9.324688478e-8   k2 = 1.193300933e-01 lk2 = -4.534370654e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.256573838e+00 ldsub = -1.405447339e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.168625007e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.510322963e-8   nfactor = {-3.309368477e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.657472975e-7   eta0 = -5.657365429e-01 leta0 = 3.143719492e-07 weta0 = 1.221245327e-21   etab = -2.105571285e-03 letab = 6.056048965e-10   u0 = 8.566582403e-03 lu0 = -1.004812388e-09 wu0 = -5.551115123e-23   ua = -4.263835804e-11 lua = -2.414708120e-16   ub = -4.555137908e-19 lub = 3.064962997e-25 wub = 1.540743956e-39 pub = 3.851859889e-46   uc = -1.047224078e-10 luc = 3.088897736e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 7.308640433e+04 lvsat = 1.651694765e-2   a0 = 1.709322966e+00 la0 = -3.259387052e-7   ags = 9.445453887e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.302213431e-01 la2 = 1.982587731e-7   b0 = 0.0   b1 = 0.0   keta = -5.758664874e-02 lketa = 7.699332989e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.886944236e-01 lpclm = 1.335541054e-7   pdiblc1 = -3.288573449e-01 lpdiblc1 = 2.184141345e-07 wpdiblc1 = 8.881784197e-22   pdiblc2 = -8.454648802e-03 lpdiblc2 = 5.071453852e-09 wpdiblc2 = -2.081668171e-23 ppdiblc2 = 6.938893904e-30   pdiblcb = -1.499370544e-01 lpdiblcb = -4.111760503e-8   drout = 4.920763650e-01 ldrout = 1.090000218e-8   pscbe1 = -6.498525204e+08 lpscbe1 = 4.317218824e+02 wpscbe1 = 1.907348633e-12 ppscbe1 = 4.768371582e-19   pscbe2 = 1.607539826e-07 lpscbe2 = -4.523478106e-14 ppscbe2 = 2.117582368e-34   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.884893411e+00 lbeta0 = 3.052351237e-7   agidl = 2.002834514e-09 lagidl = -5.967666890e-16   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.376593712e-01 lkt1 = -2.531850494e-8   kt2 = -6.756107230e-02 lkt2 = 4.391551781e-9   at = 9.442696505e+04 lat = -7.902730780e-3   ute = 4.712818972e-01 lute = -3.888555562e-07 pute = -8.881784197e-28   ua1 = 3.298078539e-09 lua1 = -8.942309315e-16   ub1 = -1.696777904e-18 lub1 = 4.548383451e-25   uc1 = -3.097635966e-11 luc1 = -1.992402306e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.160 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.078440484e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.030169421e-10   k1 = -1.029038416e+00 lk1 = 4.784953380e-7   k2 = 5.391194458e-01 lk2 = -1.703464810e-07 wk2 = 8.881784197e-22   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.925446141e+00 ldsub = -3.397181839e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.650673151e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.074904104e-8   nfactor = {4.738371709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.437660579e-7   eta0 = 4.900000008e-01 leta0 = -8.645884009e-17   etab = 2.466001640e-03 letab = -7.556952310e-10 wetab = 5.204170428e-24 petab = -4.336808690e-31   u0 = 1.371637263e-02 lu0 = -2.538291171e-9   ua = 3.518959235e-09 lua = -1.302025535e-15 pua = -3.308722450e-36   ub = -3.222538750e-18 lub = 1.130447157e-24 pub = -3.081487911e-45   uc = 3.917214497e-11 luc = -1.195922309e-17 puc = -1.938704561e-38   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.147794778e+05 lvsat = -5.545320730e-2   a0 = -2.390484591e-01 la0 = 2.542375959e-7   ags = 2.340909298e+00 lags = -2.484818634e-7   a1 = 0.0   a2 = 9.500241430e-01 la2 = -4.585800563e-8   b0 = 0.0   b1 = 0.0   keta = -9.412270452e-02 lketa = 1.857885700e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.906606977e-01 lpclm = -1.591890189e-8   pdiblc1 = 5.658853163e-01 lpdiblc1 = -4.801786142e-8   pdiblc2 = 3.245835548e-02 lpdiblc2 = -7.111415999e-9   pdiblcb = 2.481212150e+00 lpdiblcb = -8.246080592e-07 ppdiblcb = -1.776356839e-27   drout = -1.004956630e+00 ldrout = 4.566790024e-7   pscbe1 = 7.998864011e+08 lpscbe1 = 2.587501006e-2   pscbe2 = 2.085222168e-08 lpscbe2 = -3.575534212e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.071913202e+01 lbeta0 = -5.387302792e-7   agidl = -3.374235138e-09 lagidl = 1.004390227e-15 wagidl = -4.523643975e-30 pagidl = -1.815919938e-36   bgidl = 2.023190692e+09 lbgidl = -2.330572500e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.144171377e-01 lkt1 = -6.201696101e-8   kt2 = -5.940939655e-02 lkt2 = 1.964186534e-9   at = 2.293075782e+05 lat = -4.806680536e-2   ute = -1.977818730e+00 lute = 3.404253830e-7   ua1 = 1.162523927e-10 lua1 = 5.323734908e-17   ub1 = -3.497561515e-19 lub1 = 5.372894288e-26   uc1 = -3.210567629e-10 luc1 = 6.645466902e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.161 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.3e-07 wmax = 6.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-3.072770979e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.890251969e-07 wvth0 = 1.151228541e-06 pvth0 = -2.817919661e-13   k1 = 2.310038074e-01 lk1 = 2.057810293e-07 wk1 = 4.844349144e-07 pk1 = -1.185775562e-13   k2 = -1.024325072e+01 lk2 = 2.456194357e-06 wk2 = 5.782199009e-06 pk2 = -1.415337762e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.402884186e+00 ldsub = 1.428718986e-06 wdsub = 3.363389092e-06 pdsub = -8.232735649e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-3.378283995e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.217239001e-06 wvoff = 1.934444311e-05 pvoff = -4.735036061e-12   nfactor = {3.091630486e+02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.531482736e-05 wnfactor = -1.773008429e-04 pnfactor = 4.339881381e-11   eta0 = -1.144224043e+01 leta0 = 2.920714151e-06 weta0 = 6.875738768e-06 peta0 = -1.683008957e-12   etab = -6.783980956e-01 letab = 1.658464128e-07 wetab = 3.904238584e-07 petab = -9.556599995e-14   u0 = -7.026420815e-02 lu0 = 1.782860998e-08 wu0 = 4.197085066e-08 pu0 = -1.027341497e-14   ua = -6.661868955e-08 lua = 1.576874070e-14 wua = 3.712165436e-14 pua = -9.086452947e-21   ub = 1.248527572e-16 lub = -3.013481241e-23 wub = -7.094124488e-23 pub = 1.736464321e-29   uc = 5.093374037e-10 luc = -1.279365016e-16 wuc = -3.011790614e-16 puc = 7.372110475e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.768952614e+07 lvsat = -9.207995575e+00 wvsat = -2.167681219e+01 pvsat = 5.305941703e-6   a0 = 6.203842909e+00 la0 = -1.303846101e-06 wa0 = -3.069421455e-06 pa0 = 7.513176366e-13   ags = 1.250000074e+00 lags = -1.608914602e-14 wags = -2.525098353e-15 pags = 6.180869150e-22   a1 = 0.0   a2 = 8.892239722e+00 la2 = -1.993336439e-06 wa2 = -4.692571687e-06 pa2 = 1.148624235e-12   b0 = -1.461498221e-05 lb0 = 3.577382270e-12 wb0 = 8.421620427e-12 pb0 = -2.061402140e-18   b1 = 0.0   keta = 2.085331157e+00 lketa = -5.135103279e-07 wketa = -1.208869694e-06 pketa = 2.959010794e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.652099382e-01 lpclm = -1.087730038e-08 wpclm = -2.560655742e-08 ppclm = 6.267845093e-15   pdiblc1 = -6.811897704e+00 lpdiblc1 = 1.754295162e-06 wpdiblc1 = 4.129837901e-06 ppdiblc1 = -1.010881072e-12   pdiblc2 = 3.570852836e-02 lpdiblc2 = -8.437738000e-09 wpdiblc2 = -1.986353078e-08 ppdiblc2 = 4.862095747e-15   pdiblcb = 4.051562648e+01 lpdiblcb = -1.019602650e-05 wpdiblcb = -2.400276476e-05 ppdiblcb = 5.875276744e-12   drout = 1.000000068e+00 ldrout = -1.019910201e-14 wdrout = 8.282074759e-14 pdrout = -2.027245216e-20   pscbe1 = 4.669168099e+07 lpscbe1 = 1.843910438e+02 wpscbe1 = 4.340803595e+02 ppscbe1 = -1.062520200e-4   pscbe2 = 1.629049531e-07 lpscbe2 = -3.861335174e-14 wpscbe2 = -9.090082537e-14 ppscbe2 = 2.225024953e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -5.799609192e+00 lbeta0 = 3.464436437e-06 wbeta0 = 8.155730739e-06 pbeta0 = -1.996318992e-12   agidl = -4.186643252e-07 lagidl = 1.027319847e-13 wagidl = 2.418443743e-13 pagidl = -5.919745673e-20   bgidl = 1.000000468e+09 lbgidl = -1.037591705e-04 wbgidl = -6.426528931e-05 pbgidl = 1.573053741e-11   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -2.062685903e-02 lkt1 = -1.385581159e-07 wkt1 = -3.261838983e-07 pkt1 = 7.984166370e-14   kt2 = -1.709790677e+00 lkt2 = 4.060828617e-07 wkt2 = 9.559714260e-07 pkt2 = -2.339979058e-13   at = 1.485308248e+06 lat = -3.590918382e-01 wat = -8.453485956e-01 pat = 2.069202025e-7   ute = 1.204569751e+01 lute = -3.066773138e-06 wute = -7.219580679e-06 pute = 1.767172861e-12   ua1 = 1.575817723e-08 lua1 = -3.771541431e-15 wua1 = -8.878695413e-15 pua1 = 2.173282670e-21   ub1 = -2.099989256e-17 lub1 = 5.112376144e-24 wub1 = 1.203519403e-23 pub1 = -2.945914618e-30   uc1 = -5.027038166e-10 luc1 = 1.158771746e-16 wuc1 = 2.727898543e-16 puc1 = -6.677213658e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.162 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.163 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124300389e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.583094798e-7   k1 = 4.169979224e-01 lk1 = 2.938540225e-7   k2 = 5.787523347e-02 lk2 = -3.323321159e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 1.058791184e-27 pcit = -1.185846126e-32   voff = {-1.544415308e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.787950865e-7   nfactor = {1.810230600e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.882834906e-6   eta0 = 0.08   etab = -0.07   u0 = 6.082762501e-03 lu0 = 3.565351435e-8   ua = -6.616112197e-10 lua = -1.158519626e-15   ub = 4.662300295e-20 lub = 1.125904990e-23   uc = -1.046504257e-10 luc = -2.029966214e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.296000734e+04 lvsat = -2.566918583e-1   a0 = 1.627020626e+00 la0 = -3.268200833e-6   ags = 1.127420605e-01 lags = 1.098496716e-8   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 1.250763844e-07 lb0 = -1.957753127e-12 wb0 = -2.646977960e-29 pb0 = 2.117582368e-34   b1 = -6.804545270e-09 lb1 = 5.623491643e-14   keta = 3.424649349e-02 lketa = -2.182247320e-7   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 wpclm = 1.387778781e-23 ppclm = 1.110223025e-28   pdiblc1 = 0.39   pdiblc2 = 1.911548633e-03 lpdiblc2 = -1.271810464e-8   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.857143290e-09 lpscbe2 = 2.412713055e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.810749375e+01 lbeta0 = -3.630149605e-4   agidl = 2.814705940e-09 lagidl = -1.833265859e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.444100755e-01 lkt1 = 1.234958073e-7   kt2 = -6.524363936e-02 lkt2 = 1.342727668e-7   at = 7.717891133e+04 lat = -1.240739019e-1   ute = 5.643158221e-01 lute = -1.297684100e-05 wute = 5.551115123e-23   ua1 = 3.780637815e-09 lua1 = -3.388951696e-14   ub1 = -2.653212355e-18 lub1 = 2.855429361e-23   uc1 = -9.464587252e-11 luc1 = 1.300235988e-15 wuc1 = 2.584939414e-32   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.164 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140859468e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.504573657e-8   k1 = 4.604519148e-01 lk1 = -5.585393079e-8   k2 = 1.358353148e-02 lk2 = 2.411753606e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.414495418e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.214258093e-7   nfactor = {9.948645590e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.679047535e-6   eta0 = 0.08   etab = -0.07   u0 = 9.506801114e-03 lu0 = 8.097621998e-9   ua = -9.746330556e-10 lua = 1.360609680e-15   ub = 1.472299687e-18 lub = -2.144752731e-25   uc = -1.070061023e-10 luc = -1.341706802e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.345534345e+04 lvsat = -1.924496188e-2   a0 = 1.168891106e+00 la0 = 4.187224649e-7   ags = 4.434987157e-02 lags = 5.613899157e-7   a1 = 0.0   a2 = 0.8   b0 = -8.806443456e-08 lb0 = -2.424437724e-13   b1 = 3.575823691e-09 lb1 = -2.730395738e-14 wb1 = -8.271806126e-31 pb1 = 4.135903063e-36   keta = 7.542872474e-03 lketa = -3.319998307e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -4.142606150e-01 lpclm = 4.468282376e-06 wpclm = 1.110223025e-22   pdiblc1 = 0.39   pdiblc2 = 2.312663529e-04 lpdiblc2 = 8.044290883e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.465165627e-08 lpscbe2 = -2.250580619e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.011943750e-10 lalpha0 = -8.143895613e-16   alpha1 = 2.011943750e-10 lalpha1 = -8.143895613e-16   beta0 = -2.432248125e+01 lbeta0 = 2.198851815e-04 wbeta0 = 3.552713679e-21 pbeta0 = -1.421085472e-26   agidl = 6.955865393e-10 lagidl = -1.278462449e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.136981111e-01 lkt1 = -1.236671723e-7   kt2 = -3.845308193e-02 lkt2 = -8.133161144e-8   at = 2.206495351e+04 lat = 3.194708301e-1   ute = -1.923673091e+00 lute = 7.045933977e-6   ua1 = -2.981113444e-09 lua1 = 2.052753578e-14   ub1 = 2.942842689e-18 lub1 = -1.648149826e-23 wub1 = -7.703719778e-40   uc1 = 5.577709848e-10 luc1 = -3.950268087e-15 wuc1 = 2.067951531e-31 puc1 = -4.135903063e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.165 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.145429258e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.548256636e-9   k1 = 3.846063128e-01 lk1 = 2.511520008e-7   k2 = 4.228702503e-02 lk2 = -9.206774752e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.671662398e-01 ldsub = -1.243339826e-06 pdsub = -8.881784197e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.160605222e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.865677060e-8   nfactor = {2.216222452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.647344113e-7   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411601813e-01 letab = 2.880404027e-7   u0 = 1.273220293e-02 lu0 = -4.958078823e-9   ua = -3.083681764e-10 lua = -1.336280642e-15   ub = 1.131103764e-18 lub = 1.166609054e-24   uc = -1.341261632e-10 luc = 1.084341980e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.419147855e+04 lvsat = -1.031801711e-1   a0 = 1.402304588e+00 la0 = -5.260827937e-7   ags = -4.704625846e-02 lags = 9.313408859e-7   a1 = 0.0   a2 = 0.8   b0 = -1.959803238e-07 lb0 = 1.943754660e-13   b1 = -3.047654999e-09 lb1 = -4.936059274e-16   keta = 2.300377997e-02 lketa = -6.590227314e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.049877559e-01 lpclm = 3.425943017e-7   pdiblc1 = 0.39   pdiblc2 = 4.184058358e-04 lpdiblc2 = 4.693056786e-11   pdiblcb = -4.297775000e-01 lpdiblcb = 8.288932451e-7   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.707934004e-09 lpscbe2 = 1.553044224e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.023887500e-10 lalpha0 = 4.144466225e-16   alpha1 = -1.023887500e-10 lalpha1 = 4.144466225e-16   beta0 = 5.501572660e+01 lbeta0 = -1.012580327e-4   agidl = -7.892498222e-11 lagidl = 1.856585925e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.354240897e-01 lkt1 = -3.572529886e-8   kt2 = -6.326714526e-02 lkt2 = 1.911013376e-8   at = 1.633938954e+05 lat = -2.525969275e-01 wat = -1.164153218e-16   ute = -9.045128662e-02 lute = -3.745354128e-7   ua1 = 2.896511406e-09 lua1 = -3.263767152e-15 wua1 = -1.654361225e-30   ub1 = -1.914119324e-18 lub1 = 3.178391148e-24   uc1 = -8.826429466e-10 luc1 = 1.880203415e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.166 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.156253754e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.561787663e-8   k1 = 5.064465886e-01 lk1 = 1.650529987e-9   k2 = -2.574283335e-03 lk2 = -2.018817928e-10   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.600000205e-01 ldsub = -2.145607425e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.095058695e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.234316656e-9   nfactor = {2.507545012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.612974670e-7   eta0 = -5.123858625e-01 leta0 = 1.050274847e-06 weta0 = 9.194034423e-23 peta0 = 2.133709875e-28   etab = 2.826599494e-04 letab = -1.602711478e-9   u0 = 1.299327309e-02 lu0 = -5.492691778e-9   ua = -3.839322797e-10 lua = -1.181542360e-15   ub = 1.453484210e-18 lub = 5.064464363e-25   uc = -1.205586833e-10 luc = 8.065105179e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.493717597e+04 lvsat = 3.863705835e-2   a0 = 1.028226064e+00 la0 = 2.399458559e-7   ags = 2.437725462e-01 lags = 3.358094083e-7   a1 = 0.0   a2 = 0.8   b0 = -6.697383500e-09 lb0 = -1.932334070e-13   b1 = -6.829548739e-09 lb1 = 7.250861527e-15   keta = -1.770930147e-02 lketa = 1.746895719e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.234158669e-01 lpclm = -3.094748232e-7   pdiblc1 = 3.959313076e-01 lpdiblc1 = -1.214598339e-8   pdiblc2 = 4.531883283e-04 lpdiblc2 = -2.429615072e-11   pdiblcb = 1.845550000e-01 lpdiblcb = -4.291214901e-07 wpdiblcb = -2.775557562e-23   drout = 3.752086697e-01 ldrout = 3.784110665e-7   pscbe1 = 800000000.0   pscbe2 = 9.776711087e-09 lpscbe2 = -6.355707662e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.621328974e+00 lbeta0 = 1.938354859e-6   agidl = 4.019000103e-10 lagidl = 8.719645261e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.254238063e-01 lkt1 = -5.620362931e-8   kt2 = -5.956764875e-02 lkt2 = 1.153439730e-8   at = 2.776234628e+04 lat = 2.514596790e-2   ute = 5.384763382e-01 lute = -1.662437680e-6   ua1 = 3.118603033e-09 lua1 = -3.718560834e-15   ub1 = -1.637022257e-18 lub1 = 2.610958703e-24 pub1 = 7.703719778e-46   uc1 = 2.633427840e-12 luc1 = 6.735658696e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.167 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.189894012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.086529730e-8   k1 = 5.880791324e-01 lk1 = -8.388200862e-8   k2 = -4.584297371e-02 lk2 = 4.513397027e-08 wk2 = -6.938893904e-24 pk2 = -8.673617380e-30   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.507070000e-01 ldsub = 8.494385269e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.503262196e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.800485898e-8   nfactor = {2.363154285e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.100084730e-7   eta0 = 1.017868271e+00 leta0 = -5.530871778e-7   etab = -1.517546071e-03 letab = 2.834993852e-10   u0 = 8.867175292e-03 lu0 = -1.169469657e-9   ua = -2.637979932e-09 lua = 1.180192418e-15   ub = 3.944787243e-18 lub = -2.103878599e-24   uc = -3.838396610e-11 luc = -5.449562538e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.527989752e+03 lvsat = 5.903217237e-2   a0 = 1.413819476e+00 la0 = -1.640692811e-7   ags = -1.869811243e-01 lags = 7.871423354e-7   a1 = 0.0   a2 = 1.137258461e+00 la2 = -3.533709843e-7   b0 = -4.005015160e-07 lb0 = 2.193847179e-13   b1 = 1.900621939e-10 lb1 = -1.041113183e-16   keta = 4.551757475e-02 lketa = -4.877858303e-08 wketa = 6.071532166e-24 pketa = 1.040834086e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 8.422820869e-01 lpclm = -2.244648769e-7   pdiblc1 = 7.288532800e-01 lpdiblc1 = -3.609733030e-7   pdiblc2 = 2.066929197e-05 lpdiblc2 = 4.288864826e-10   pdiblcb = -0.225   drout = 9.821963946e-01 ldrout = -2.575754971e-7   pscbe1 = 1.524942164e+09 lpscbe1 = -7.595762759e+2   pscbe2 = -6.642801811e-08 lpscbe2 = 7.920983936e-14 wpscbe2 = 1.323488980e-29 ppscbe2 = -1.323488980e-35   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.312170425e+00 lbeta0 = 2.262283457e-6   agidl = 1.585458645e-09 lagidl = -3.681386223e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.737893819e-01 lkt1 = -5.527388326e-9   kt2 = -3.652476254e-02 lkt2 = -1.260936280e-8   at = 2.082532054e+04 lat = 3.241441004e-2   ute = -1.935073039e+00 lute = 9.292855189e-7   ua1 = -2.726681161e-09 lua1 = 2.405981813e-15 wua1 = -8.271806126e-31 pua1 = -4.135903063e-37   ub1 = 2.740683756e-18 lub1 = -1.975892216e-24   uc1 = 2.140158506e-10 luc1 = -1.541246310e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.168 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.122397186e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.389222392e-8   k1 = 2.647184581e-01 lk1 = 9.324688478e-8   k2 = 1.193300933e-01 lk2 = -4.534370654e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.256573838e+00 ldsub = -1.405447339e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.168625007e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.510322963e-8   nfactor = {-3.309368477e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.657472975e-7   eta0 = -5.657365429e-01 leta0 = 3.143719492e-07 weta0 = -9.020562075e-23 peta0 = 7.285838599e-29   etab = -2.105571285e-03 letab = 6.056048965e-10 petab = -4.336808690e-31   u0 = 8.566582403e-03 lu0 = -1.004812388e-9   ua = -4.263835804e-11 lua = -2.414708120e-16   ub = -4.555137908e-19 lub = 3.064962997e-25 pub = 4.814824861e-47   uc = -1.047224078e-10 luc = 3.088897736e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 7.308640433e+04 lvsat = 1.651694765e-2   a0 = 1.709322966e+00 la0 = -3.259387052e-7   ags = 9.445453887e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.302213431e-01 la2 = 1.982587731e-7   b0 = 0.0   b1 = 0.0   keta = -5.758664874e-02 lketa = 7.699332989e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.886944236e-01 lpclm = 1.335541054e-7   pdiblc1 = -3.288573449e-01 lpdiblc1 = 2.184141345e-07 ppdiblc1 = 5.551115123e-29   pdiblc2 = -8.454648802e-03 lpdiblc2 = 5.071453852e-09 wpdiblc2 = -1.734723476e-24 ppdiblc2 = -1.517883041e-30   pdiblcb = -1.499370544e-01 lpdiblcb = -4.111760503e-8   drout = 4.920763650e-01 ldrout = 1.090000218e-8   pscbe1 = -6.498525204e+08 lpscbe1 = 4.317218824e+02 ppscbe1 = -5.960464478e-20   pscbe2 = 1.607539826e-07 lpscbe2 = -4.523478106e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.884893411e+00 lbeta0 = 3.052351237e-7   agidl = 2.002834514e-09 lagidl = -5.967666890e-16   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.376593712e-01 lkt1 = -2.531850494e-8   kt2 = -6.756107230e-02 lkt2 = 4.391551781e-9   at = 9.442696505e+04 lat = -7.902730780e-3   ute = 4.712818972e-01 lute = -3.888555562e-7   ua1 = 3.298078539e-09 lua1 = -8.942309315e-16   ub1 = -1.696777904e-18 lub1 = 4.548383451e-25   uc1 = -3.097635966e-11 luc1 = -1.992402306e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.169 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.078440484e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.030169421e-10   k1 = -1.029038416e+00 lk1 = 4.784953380e-7   k2 = 5.391194458e-01 lk2 = -1.703464810e-07 wk2 = 1.110223025e-22   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.925446141e+00 ldsub = -3.397181839e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.650673151e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.074904104e-8   nfactor = {4.738371709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.437660579e-7   eta0 = 4.900000008e-01 leta0 = -8.645972827e-17   etab = 2.466001640e-03 letab = -7.556952310e-10 wetab = -4.336808690e-25 petab = 5.421010862e-32   u0 = 1.371637263e-02 lu0 = -2.538291171e-9   ua = 3.518959235e-09 lua = -1.302025535e-15 pua = -4.135903063e-37   ub = -3.222538750e-18 lub = 1.130447157e-24   uc = 3.917214497e-11 luc = -1.195922309e-17 wuc = 4.846761402e-33 puc = 3.231174268e-39   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.147794778e+05 lvsat = -5.545320730e-2   a0 = -2.390484591e-01 la0 = 2.542375959e-7   ags = 2.340909298e+00 lags = -2.484818634e-7   a1 = 0.0   a2 = 9.500241430e-01 la2 = -4.585800563e-8   b0 = 0.0   b1 = 0.0   keta = -9.412270452e-02 lketa = 1.857885700e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.906606977e-01 lpclm = -1.591890189e-8   pdiblc1 = 5.658853163e-01 lpdiblc1 = -4.801786142e-8   pdiblc2 = 3.245835548e-02 lpdiblc2 = -7.111415999e-09 ppdiblc2 = 3.469446952e-30   pdiblcb = 2.481212150e+00 lpdiblcb = -8.246080592e-07 wpdiblcb = 8.881784197e-22 ppdiblcb = 1.110223025e-28   drout = -1.004956630e+00 ldrout = 4.566790024e-7   pscbe1 = 7.998864011e+08 lpscbe1 = 2.587501006e-2   pscbe2 = 2.085222168e-08 lpscbe2 = -3.575534212e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.071913202e+01 lbeta0 = -5.387302792e-7   agidl = -3.374235138e-09 lagidl = 1.004390227e-15 wagidl = 4.426708747e-31 pagidl = 4.846761402e-38   bgidl = 2.023190692e+09 lbgidl = -2.330572500e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.144171377e-01 lkt1 = -6.201696101e-8   kt2 = -5.940939655e-02 lkt2 = 1.964186534e-9   at = 2.293075782e+05 lat = -4.806680536e-2   ute = -1.977818730e+00 lute = 3.404253830e-7   ua1 = 1.162523927e-10 lua1 = 5.323734908e-17   ub1 = -3.497561515e-19 lub1 = 5.372894288e-26   uc1 = -3.210567629e-10 luc1 = 6.645466902e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.170 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.3e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {1.093740355e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.898843489e-07 wvth0 = -6.506037946e-07 pvth0 = 1.592515438e-13   k1 = 2.423321921e-01 lk1 = 2.030081240e-07 wk1 = 4.780204205e-07 pk1 = -1.170074484e-13   k2 = 1.262345327e+00 lk2 = -3.600879153e-07 wk2 = -7.326376512e-07 pk2 = 1.793313811e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.324232323e+00 ldsub = 1.409466976e-06 wdsub = 3.318853890e-06 pdsub = -8.123724609e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {4.222291933e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.085467156e-06 wvoff = -2.175278731e-06 pvoff = 5.324538513e-13   nfactor = {-3.769143814e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.586479627e-06 wnfactor = 1.909926685e-05 pnfactor = -4.675023043e-12   eta0 = -1.128145435e+01 leta0 = 2.881357739e-06 weta0 = 6.784696546e-06 peta0 = -1.660724097e-12   etab = -6.692680777e-01 letab = 1.636116127e-07 wetab = 3.852541502e-07 petab = -9.430058461e-14   u0 = -3.150663768e-02 lu0 = 8.341725670e-09 wu0 = 2.002507401e-08 pu0 = -4.901637492e-15   ua = -1.532665298e-08 lua = 3.213732445e-15 wua = 8.078461909e-15 pua = -1.977405514e-21   ub = 1.144422675e-17 lub = -2.375239382e-24 wub = -6.725705884e-24 pub = 1.646284658e-30   uc = 5.022944134e-10 luc = -1.262125536e-16 wuc = -2.971910949e-16 puc = 7.274495025e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -9.773385109e+05 lvsat = 2.566862201e-01 wvsat = 2.176039206e-01 pvsat = -5.326399966e-8   a0 = 6.132065760e+00 la0 = -1.286276850e-06 wa0 = -3.028778936e-06 pa0 = 7.413693642e-13   ags = 1.250000069e+00 lags = -1.488242241e-14 wags = 2.663398391e-16 pags = -6.519318418e-23   a1 = 0.0   a2 = 8.782505590e+00 la2 = -1.966476267e-06 wa2 = -4.630436710e-06 pa2 = 1.133415146e-12   b0 = 1.826872776e-06 lb0 = -4.471727837e-13 wb0 = -8.882840036e-13 pb0 = 2.174297170e-19   b1 = 0.0   keta = 2.057061952e+00 lketa = -5.065907333e-07 wketa = -1.192862766e-06 pketa = 2.919829835e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.646111422e-01 lpclm = -1.073073008e-08 wpclm = -2.526749994e-08 ppclm = 6.184852299e-15   pdiblc1 = -6.715322679e+00 lpdiblc1 = 1.730656010e-06 wpdiblc1 = 4.075154032e-06 ppdiblc1 = -9.974958281e-13   pdiblc2 = 3.524401915e-02 lpdiblc2 = -8.324037759e-09 wpdiblc2 = -1.960051080e-08 ppdiblc2 = 4.797715032e-15   pdiblcb = 3.995433271e+01 lpdiblcb = -1.005863581e-05 wpdiblcb = -2.368494226e-05 ppdiblcb = 5.797481743e-12   drout = 1.000000229e+00 ldrout = -4.977779788e-14 wdrout = -8.735650425e-15 pdrout = 2.138269117e-21   pscbe1 = 5.684258016e+07 lpscbe1 = 1.819063575e+02 wpscbe1 = 4.283325956e+02 ppscbe1 = -1.048451111e-4   pscbe2 = 1.607792351e-07 lpscbe2 = -3.809302913e-14 wpscbe2 = -8.969717584e-14 ppscbe2 = 2.195562622e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = -5.608890329e+00 lbeta0 = 3.417753227e-06 wbeta0 = 8.047739616e-06 pbeta0 = -1.969885464e-12   agidl = 5.499990701e-08 lagidl = -1.320917770e-14 wagidl = -2.635947117e-14 pagidl = 6.452139555e-21   bgidl = 1.000000342e+09 lbgidl = -7.304783249e-05 wbgidl = 6.778484344e-06 pbgidl = -1.659203529e-12   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -2.825465909e-02 lkt1 = -1.366910211e-07 wkt1 = -3.218647938e-07 pkt1 = 7.878445490e-14   kt2 = -1.687435397e+00 lkt2 = 4.006108479e-07 wkt2 = 9.433131508e-07 pkt2 = -2.308994765e-13   at = 1.465539918e+06 lat = -3.542530451e-01 wat = -8.341551343e-01 pat = 2.041803230e-7   ute = 1.187687052e+01 lute = -3.025448511e-06 wute = -7.123985433e-06 pute = 1.743773534e-12   ua1 = 1.555055545e-08 lua1 = -3.720720810e-15 wua1 = -8.761133317e-15 pua1 = 2.144506408e-21   ub1 = -2.071844854e-17 lub1 = 5.043485685e-24 wub1 = 1.187583142e-23 pub1 = -2.906906636e-30   uc1 = -4.963247131e-10 luc1 = 1.143157295e-16 wuc1 = 2.691778018e-16 puc1 = -6.588799643e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.171 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.172 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.124300389e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.583094798e-7   k1 = 4.169979224e-01 lk1 = 2.938540225e-7   k2 = 5.787523347e-02 lk2 = -3.323321159e-07 wk2 = 2.220446049e-22   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = 1.016439537e-26 pcit = 1.897353802e-31   voff = {-1.544415308e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.787950865e-7   nfactor = {1.810230600e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.882834906e-6   eta0 = 0.08   etab = -0.07   u0 = 6.082762501e-03 lu0 = 3.565351435e-8   ua = -6.616112197e-10 lua = -1.158519626e-15   ub = 4.662300295e-20 lub = 1.125904990e-23 pub = -2.465190329e-44   uc = -1.046504257e-10 luc = -2.029966214e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.296000734e+04 lvsat = -2.566918583e-1   a0 = 1.627020626e+00 la0 = -3.268200833e-6   ags = 1.127420605e-01 lags = 1.098496716e-8   a1 = 0.0   a2 = 1.084010146e+00 la2 = -2.285649751e-6   b0 = 1.250763844e-07 lb0 = -1.957753127e-12 wb0 = -2.117582368e-28 pb0 = 1.694065895e-33   b1 = -6.804545270e-09 lb1 = 5.623491643e-14   keta = 3.424649349e-02 lketa = -2.182247320e-07 pketa = 8.881784197e-28   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -6.947412752e-02 lpclm = 1.693518302e-06 ppclm = 2.664535259e-27   pdiblc1 = 0.39   pdiblc2 = 1.911548633e-03 lpdiblc2 = -1.271810464e-08 wpdiblc2 = -6.938893904e-24   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.857143290e-09 lpscbe2 = 2.412713055e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -6.706479167e-11 lalpha0 = 1.344499854e-15   alpha1 = -6.706479167e-11 lalpha1 = 1.344499854e-15   beta0 = 4.810749375e+01 lbeta0 = -3.630149605e-4   agidl = 2.814705940e-09 lagidl = -1.833265859e-14 wagidl = 1.323488980e-29   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.444100755e-01 lkt1 = 1.234958073e-7   kt2 = -6.524363936e-02 lkt2 = 1.342727668e-7   at = 7.717891133e+04 lat = -1.240739019e-1   ute = 5.643158221e-01 lute = -1.297684100e-05 wute = 4.440892099e-22 pute = 1.421085472e-26   ua1 = 3.780637815e-09 lua1 = -3.388951696e-14   ub1 = -2.653212355e-18 lub1 = 2.855429361e-23 wub1 = 6.162975822e-39 pub1 = -4.930380658e-44   uc1 = -9.464587252e-11 luc1 = 1.300235988e-15 wuc1 = 2.067951531e-31 puc1 = -3.308722450e-36   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.173 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.140859468e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.504573657e-8   k1 = 4.604519148e-01 lk1 = -5.585393079e-8   k2 = 1.358353148e-02 lk2 = 2.411753606e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.414495418e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.214258093e-7   nfactor = {9.948645590e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.679047535e-6   eta0 = 0.08   etab = -0.07   u0 = 9.506801114e-03 lu0 = 8.097621998e-9   ua = -9.746330556e-10 lua = 1.360609680e-15   ub = 1.472299687e-18 lub = -2.144752731e-25   uc = -1.070061023e-10 luc = -1.341706802e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.345534345e+04 lvsat = -1.924496188e-2   a0 = 1.168891106e+00 la0 = 4.187224649e-7   ags = 4.434987157e-02 lags = 5.613899157e-7   a1 = 0.0   a2 = 0.8   b0 = -8.806443456e-08 lb0 = -2.424437724e-13   b1 = 3.575823691e-09 lb1 = -2.730395738e-14 wb1 = -3.308722450e-30 pb1 = -5.293955920e-35   keta = 7.542872474e-03 lketa = -3.319998307e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -4.142606150e-01 lpclm = 4.468282376e-06 ppclm = 3.552713679e-27   pdiblc1 = 0.39   pdiblc2 = 2.312663529e-04 lpdiblc2 = 8.044290883e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.465165627e-08 lpscbe2 = -2.250580619e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.011943750e-10 lalpha0 = -8.143895613e-16   alpha1 = 2.011943750e-10 lalpha1 = -8.143895613e-16   beta0 = -2.432248125e+01 lbeta0 = 2.198851815e-04 wbeta0 = -5.684341886e-20 pbeta0 = 1.136868377e-25   agidl = 6.955865393e-10 lagidl = -1.278462449e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.136981111e-01 lkt1 = -1.236671723e-7   kt2 = -3.845308193e-02 lkt2 = -8.133161144e-8   at = 2.206495351e+04 lat = 3.194708301e-1   ute = -1.923673091e+00 lute = 7.045933977e-6   ua1 = -2.981113444e-09 lua1 = 2.052753578e-14 wua1 = -3.308722450e-30 pua1 = -2.646977960e-35   ub1 = 2.942842689e-18 lub1 = -1.648149826e-23 pub1 = -2.465190329e-44   uc1 = 5.577709848e-10 luc1 = -3.950268087e-15 wuc1 = 4.135903063e-31 puc1 = 4.963083675e-36   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.174 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.145429258e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.548256636e-9   k1 = 3.846063128e-01 lk1 = 2.511520008e-7   k2 = 4.228702503e-02 lk2 = -9.206774752e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.671662398e-01 ldsub = -1.243339826e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.160605222e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.865677060e-8   nfactor = {2.216222452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.647344113e-7   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411601813e-01 letab = 2.880404027e-7   u0 = 1.273220293e-02 lu0 = -4.958078823e-9   ua = -3.083681764e-10 lua = -1.336280642e-15   ub = 1.131103764e-18 lub = 1.166609054e-24   uc = -1.341261632e-10 luc = 1.084341980e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.419147855e+04 lvsat = -1.031801711e-1   a0 = 1.402304588e+00 la0 = -5.260827937e-7   ags = -4.704625846e-02 lags = 9.313408859e-7   a1 = 0.0   a2 = 0.8   b0 = -1.959803238e-07 lb0 = 1.943754660e-13   b1 = -3.047654999e-09 lb1 = -4.936059274e-16   keta = 2.300377997e-02 lketa = -6.590227314e-08 wketa = -5.551115123e-23   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.049877559e-01 lpclm = 3.425943017e-7   pdiblc1 = 0.39   pdiblc2 = 4.184058358e-04 lpdiblc2 = 4.693056786e-11   pdiblcb = -4.297775000e-01 lpdiblcb = 8.288932451e-7   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 8.707934004e-09 lpscbe2 = 1.553044224e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.023887500e-10 lalpha0 = 4.144466225e-16   alpha1 = -1.023887500e-10 lalpha1 = 4.144466225e-16   beta0 = 5.501572660e+01 lbeta0 = -1.012580327e-4   agidl = -7.892498222e-11 lagidl = 1.856585925e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.354240898e-01 lkt1 = -3.572529886e-8   kt2 = -6.326714526e-02 lkt2 = 1.911013376e-8   at = 1.633938953e+05 lat = -2.525969275e-1   ute = -9.045128663e-02 lute = -3.745354128e-7   ua1 = 2.896511406e-09 lua1 = -3.263767152e-15   ub1 = -1.914119324e-18 lub1 = 3.178391148e-24 pub1 = -1.232595164e-44   uc1 = -8.826429466e-10 luc1 = 1.880203415e-15   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.175 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.156253754e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.561787663e-8   k1 = 5.064465886e-01 lk1 = 1.650529987e-9   k2 = -2.574283335e-03 lk2 = -2.018817928e-10   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.600000205e-01 ldsub = -2.145607425e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.095058695e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.234316656e-9   nfactor = {2.507545012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.612974670e-7   eta0 = -5.123858625e-01 leta0 = 1.050274847e-06 weta0 = 1.838806885e-22 peta0 = -1.592476151e-27   etab = 2.826599494e-04 letab = -1.602711478e-09 petab = -3.469446952e-30   u0 = 1.299327309e-02 lu0 = -5.492691778e-9   ua = -3.839322797e-10 lua = -1.181542360e-15   ub = 1.453484210e-18 lub = 5.064464363e-25   uc = -1.205586833e-10 luc = 8.065105179e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.493717597e+04 lvsat = 3.863705835e-2   a0 = 1.028226064e+00 la0 = 2.399458559e-7   ags = 2.437725462e-01 lags = 3.358094083e-7   a1 = 0.0   a2 = 0.8   b0 = -6.697383500e-09 lb0 = -1.932334070e-13   b1 = -6.829548739e-09 lb1 = 7.250861527e-15   keta = -1.770930147e-02 lketa = 1.746895719e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.234158669e-01 lpclm = -3.094748232e-7   pdiblc1 = 3.959313076e-01 lpdiblc1 = -1.214598339e-8   pdiblc2 = 4.531883283e-04 lpdiblc2 = -2.429615072e-11   pdiblcb = 1.845550000e-01 lpdiblcb = -4.291214901e-07 wpdiblcb = -2.220446049e-22 ppdiblcb = -4.440892099e-28   drout = 3.752086697e-01 ldrout = 3.784110665e-7   pscbe1 = 800000000.0   pscbe2 = 9.776711087e-09 lpscbe2 = -6.355707662e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.621328974e+00 lbeta0 = 1.938354859e-6   agidl = 4.019000103e-10 lagidl = 8.719645261e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.254238063e-01 lkt1 = -5.620362931e-8   kt2 = -5.956764875e-02 lkt2 = 1.153439730e-8   at = 2.776234628e+04 lat = 2.514596790e-2   ute = 5.384763382e-01 lute = -1.662437680e-06 pute = -3.552713679e-27   ua1 = 3.118603033e-09 lua1 = -3.718560834e-15   ub1 = -1.637022257e-18 lub1 = 2.610958703e-24 wub1 = 3.081487911e-39 pub1 = -6.162975822e-45   uc1 = 2.633427840e-12 luc1 = 6.735658696e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.176 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.189894012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.086529730e-8   k1 = 5.880791324e-01 lk1 = -8.388200862e-8   k2 = -4.584297371e-02 lk2 = 4.513397027e-08 wk2 = 2.775557562e-23 pk2 = -8.326672685e-29   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.507070000e-01 ldsub = 8.494385269e-07 pdsub = -8.881784197e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.503262196e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.800485898e-8   nfactor = {2.363154285e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.100084730e-7   eta0 = 1.017868271e+00 leta0 = -5.530871778e-7   etab = -1.517546071e-03 letab = 2.834993852e-10   u0 = 8.867175292e-03 lu0 = -1.169469657e-9   ua = -2.637979932e-09 lua = 1.180192418e-15   ub = 3.944787243e-18 lub = -2.103878599e-24   uc = -3.838396610e-11 luc = -5.449562538e-18   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -4.527989752e+03 lvsat = 5.903217237e-2   a0 = 1.413819476e+00 la0 = -1.640692811e-7   ags = -1.869811243e-01 lags = 7.871423354e-07 pags = 1.776356839e-27   a1 = 0.0   a2 = 1.137258461e+00 la2 = -3.533709843e-7   b0 = -4.005015160e-07 lb0 = 2.193847179e-13   b1 = 1.900621939e-10 lb1 = -1.041113183e-16   keta = 4.551757475e-02 lketa = -4.877858303e-08 wketa = -1.110223025e-22 pketa = 3.816391647e-29   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 8.422820869e-01 lpclm = -2.244648769e-7   pdiblc1 = 7.288532800e-01 lpdiblc1 = -3.609733030e-7   pdiblc2 = 2.066929197e-05 lpdiblc2 = 4.288864826e-10   pdiblcb = -0.225   drout = 9.821963946e-01 ldrout = -2.575754971e-7   pscbe1 = 1.524942164e+09 lpscbe1 = -7.595762759e+2   pscbe2 = -6.642801811e-08 lpscbe2 = 7.920983936e-14 wpscbe2 = -5.293955920e-29 ppscbe2 = -5.293955920e-35   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 4.312170425e+00 lbeta0 = 2.262283457e-6   agidl = 1.585458645e-09 lagidl = -3.681386223e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.737893819e-01 lkt1 = -5.527388326e-9   kt2 = -3.652476254e-02 lkt2 = -1.260936280e-8   at = 2.082532054e+04 lat = 3.241441004e-2   ute = -1.935073039e+00 lute = 9.292855189e-7   ua1 = -2.726681161e-09 lua1 = 2.405981813e-15 wua1 = -3.308722450e-30 pua1 = -3.308722450e-36   ub1 = 2.740683756e-18 lub1 = -1.975892216e-24 wub1 = -6.162975822e-39   uc1 = 2.140158506e-10 luc1 = -1.541246310e-16 wuc1 = 4.135903063e-31   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.177 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.122397186e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.389222392e-8   k1 = 2.647184581e-01 lk1 = 9.324688478e-8   k2 = 1.193300933e-01 lk2 = -4.534370654e-08 wk2 = 2.220446049e-22   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.256573838e+00 ldsub = -1.405447339e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.168625007e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.510322963e-8   nfactor = {-3.309368477e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.657472975e-7   eta0 = -5.657365429e-01 leta0 = 3.143719492e-07 weta0 = 8.881784197e-22 peta0 = -1.110223025e-28   etab = -2.105571285e-03 letab = 6.056048965e-10   u0 = 8.566582403e-03 lu0 = -1.004812388e-9   ua = -4.263835804e-11 lua = -2.414708120e-16   ub = -4.555137908e-19 lub = 3.064962997e-25 wub = 7.703719778e-40 pub = -1.925929944e-46   uc = -1.047224078e-10 luc = 3.088897736e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 7.308640433e+04 lvsat = 1.651694765e-2   a0 = 1.709322966e+00 la0 = -3.259387052e-7   ags = 9.445453887e-01 lags = 1.673203997e-7   a1 = 0.0   a2 = 1.302213431e-01 la2 = 1.982587731e-7   b0 = 0.0   b1 = 0.0   keta = -5.758664874e-02 lketa = 7.699332989e-9   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.886944236e-01 lpclm = 1.335541054e-7   pdiblc1 = -3.288573449e-01 lpdiblc1 = 2.184141345e-7   pdiblc2 = -8.454648802e-03 lpdiblc2 = 5.071453852e-09 ppdiblc2 = -3.469446952e-30   pdiblcb = -1.499370544e-01 lpdiblcb = -4.111760503e-8   drout = 4.920763650e-01 ldrout = 1.090000218e-8   pscbe1 = -6.498525204e+08 lpscbe1 = 4.317218824e+02 ppscbe1 = 2.384185791e-19   pscbe2 = 1.607539826e-07 lpscbe2 = -4.523478106e-14   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.884893411e+00 lbeta0 = 3.052351237e-7   agidl = 2.002834514e-09 lagidl = -5.967666890e-16   bgidl = 7.135065664e+08 lbgidl = 1.569339406e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.376593712e-01 lkt1 = -2.531850494e-8   kt2 = -6.756107230e-02 lkt2 = 4.391551781e-9   at = 9.442696505e+04 lat = -7.902730780e-03 wat = -4.656612873e-16   ute = 4.712818972e-01 lute = -3.888555562e-07 pute = -8.881784197e-28   ua1 = 3.298078539e-09 lua1 = -8.942309315e-16   ub1 = -1.696777904e-18 lub1 = 4.548383451e-25   uc1 = -3.097635966e-11 luc1 = -1.992402306e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.178 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.078440484e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.030169421e-10   k1 = -1.029038416e+00 lk1 = 4.784953380e-7   k2 = 5.391194458e-01 lk2 = -1.703464810e-07 pk2 = -1.110223025e-28   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.925446141e+00 ldsub = -3.397181839e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.650673151e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.074904104e-8   nfactor = {4.738371709e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.437660579e-7   eta0 = 4.900000008e-01 leta0 = -8.645884009e-17   etab = 2.466001640e-03 letab = -7.556952310e-10 wetab = 1.734723476e-24 petab = -1.301042607e-30   u0 = 1.371637263e-02 lu0 = -2.538291171e-9   ua = 3.518959235e-09 lua = -1.302025535e-15 pua = 3.308722450e-36   ub = -3.222538750e-18 lub = 1.130447157e-24   uc = 3.917214497e-11 luc = -1.195922309e-17 wuc = -3.877409121e-32 puc = -6.462348536e-39   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.147794778e+05 lvsat = -5.545320730e-2   a0 = -2.390484591e-01 la0 = 2.542375959e-7   ags = 2.340909298e+00 lags = -2.484818634e-7   a1 = 0.0   a2 = 9.500241430e-01 la2 = -4.585800563e-8   b0 = 0.0   b1 = 0.0   keta = -9.412270452e-02 lketa = 1.857885700e-08 wketa = 4.440892099e-22   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.906606977e-01 lpclm = -1.591890189e-8   pdiblc1 = 5.658853163e-01 lpdiblc1 = -4.801786142e-8   pdiblc2 = 3.245835548e-02 lpdiblc2 = -7.111415999e-09 wpdiblc2 = 1.110223025e-22   pdiblcb = 2.481212150e+00 lpdiblcb = -8.246080592e-07 wpdiblcb = 3.552713679e-21 ppdiblcb = -8.881784197e-28   drout = -1.004956630e+00 ldrout = 4.566790024e-7   pscbe1 = 7.998864011e+08 lpscbe1 = 2.587501006e-2   pscbe2 = 2.085222168e-08 lpscbe2 = -3.575534212e-15 wpscbe2 = -1.058791184e-28   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.071913202e+01 lbeta0 = -5.387302792e-7   agidl = -3.374235138e-09 lagidl = 1.004390227e-15 wagidl = -4.652890946e-31 pagidl = 6.074607623e-37   bgidl = 2.023190692e+09 lbgidl = -2.330572500e+2   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710448227029   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.70969974265993e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.144171377e-01 lkt1 = -6.201696101e-8   kt2 = -5.940939655e-02 lkt2 = 1.964186534e-9   at = 2.293075782e+05 lat = -4.806680536e-2   ute = -1.977818730e+00 lute = 3.404253830e-7   ua1 = 1.162523927e-10 lua1 = 5.323734908e-17   ub1 = -3.497561515e-19 lub1 = 5.372894288e-26   uc1 = -3.210567629e-10 luc1 = 6.645466902e-17   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.179 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.547845422e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.525626313e-06 wvth0 = 6.928697116e-06 pvth0 = -1.695971837e-12   k1 = -3.535511583e-01 lk1 = 3.488654711e-07 wk1 = 7.677579737e-07 pk1 = -1.879279580e-13   k2 = -1.138031412e+01 lk2 = 2.734519051e-06 wk2 = 5.414627937e-06 pk2 = -1.325365553e-12   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 5.579725854e+00 ldsub = -1.259549387e-06 wdsub = -1.982999502e-06 pdsub = 4.853887032e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-3.060781583e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.440072472e-06 wvoff = 1.476023423e-05 pvoff = -3.612936333e-12   nfactor = {3.152322061e+02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.680040539e-05 wnfactor = -1.525035025e-04 pnfactor = 3.732904483e-11   eta0 = 8.825881263e+00 leta0 = -2.040415336e-06 weta0 = -2.992133464e-06 peta0 = 7.323994687e-13   etab = 4.770600832e-01 letab = -1.169808629e-07 wetab = -1.721272842e-07 petab = 4.213245598e-14   u0 = 4.379060520e-01 lu0 = -1.065587654e-07 wu0 = -2.082183969e-07 pu0 = 5.096665811e-14   ua = 1.720794081e-07 lua = -4.265858615e-14 wua = -8.304436198e-14 pua = 2.032718370e-20   ub = -1.164405199e-16 lub = 2.892774947e-23 wub = 5.545595024e-23 pub = -1.357423022e-29   uc = -4.961458717e-10 luc = 1.181806672e-16 wuc = 1.882825218e-16 puc = -4.608685428e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.081509976e+07 lvsat = -7.525307859e+00 wvsat = -1.524089693e+01 pvsat = 3.730590545e-6   a0 = -2.630163620e-01 la0 = 2.790793767e-07 wa0 = 8.071463387e-08 pa0 = -1.975692451e-14   ags = 1.249999927e+00 lags = 1.989990039e-14 wags = 6.935948704e-14 pags = -1.697746654e-20   a1 = 0.0   a2 = -7.253433966e+00 la2 = 1.958720838e-06 wa2 = 3.166750253e-06 pa2 = -7.751412931e-13   b0 = -2.765724960e-05 lb0 = 6.769803270e-12 wb0 = 1.344783979e-11 pb0 = -3.291694984e-18   b1 = 0.0   keta = -1.572647300e+00 lketa = 3.818713489e-07 wketa = 5.720180234e-07 pketa = -1.400157117e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 6.664325522e-01 lpclm = -1.117656572e-08 wpclm = -2.615312779e-08 ppclm = 6.401631856e-15   pdiblc1 = 1.489156711e+00 lpdiblc1 = -2.775954329e-07 wpdiblc1 = 8.587360872e-08 ppdiblc1 = -2.101971258e-14   pdiblc2 = 2.699551403e-02 lpdiblc2 = -6.305009917e-09 wpdiblc2 = -1.558982366e-08 ppdiblc2 = 3.815999086e-15   pdiblcb = -1.746331918e+01 lpdiblcb = 3.995769929e-06 wpdiblcb = 4.233357451e-06 ppdiblcb = -1.036220070e-12   drout = 1.000000066e+00 ldrout = -9.724544725e-15 wdrout = 7.082795150e-14 pdrout = -1.733690880e-20   pscbe1 = 1.326253667e+09 lpscbe1 = -1.288137414e+02 wpscbe1 = -1.888956961e+02 ppscbe1 = 4.623694401e-5   pscbe2 = -1.789199051e-08 lpscbe2 = 5.641220131e-15 wpscbe2 = -2.821508449e-15 ppscbe2 = 6.906347306e-22   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.880698925e+01 lbeta0 = -2.558643698e-06 wbeta0 = -3.824042346e-06 pbeta0 = 9.360299652e-13   agidl = -3.639718934e-07 lagidl = 8.934464475e-14 wagidl = 1.773580253e-13 pagidl = -4.341281064e-20   bgidl = 1.000000455e+09 lbgidl = -1.007603912e-04 wbgidl = -4.827099609e-05 pbgidl = 1.181552887e-11   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 3.210489251e-01 lkt1 = -2.221918059e-07 wkt1 = -4.917073741e-07 pkt1 = 1.203576725e-13   kt2 = 1.148755897e+00 lkt2 = -2.936178759e-07 wkt2 = -4.357338142e-07 pkt2 = 1.066567444e-13   at = -6.256238753e+05 lat = 1.576115724e-01 wat = 1.826356193e-01 pat = -4.470463371e-8   ute = -2.774541501e+00 lute = 5.608508671e-07 wute = -6.286384746e-14 pute = 1.538749572e-20   ua1 = -4.447390893e-10 lua1 = 1.945274117e-16 wua1 = -9.837092617e-16 pua1 = 2.407874345e-22   ub1 = 4.067342155e-18 lub1 = -1.023456232e-24 wub1 = -1.758131610e-25 pub1 = 4.303466648e-32   uc1 = -7.784437474e-10 luc1 = 1.833714161e-16 wuc1 = 4.063531040e-16 puc1 = -9.946508104e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.180 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.181 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.130220088e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.963269289e-08 wvth0 = 2.819149934e-09 pvth0 = -5.651768358e-14   k1 = 3.731509609e-01 lk1 = 1.172888042e-06 wk1 = 2.088132619e-08 pk1 = -4.186241291e-13   k2 = 8.027333534e-02 lk2 = -7.813642227e-07 wk2 = -1.066669285e-08 pk2 = 2.138434583e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 pcit = -5.082197684e-33   voff = {-1.361852111e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.447936747e-07 wvoff = -8.694243607e-09 pvoff = 1.743002396e-13   nfactor = {1.657449059e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.180095061e-06 wnfactor = 7.275945905e-08 pnfactor = -1.458665264e-12   eta0 = 0.08   etab = -0.07   u0 = 1.472877300e-03 lu0 = 1.280714556e-07 wu0 = 2.195374849e-09 pu0 = -4.401238102e-14   ua = -2.475803199e-10 lua = -9.458917947e-15 wua = -1.971747634e-16 pua = 3.952915293e-21   ub = -1.830092570e-18 lub = 4.888302146e-23 wub = 8.937520109e-25 pub = -1.791773922e-29   uc = -1.100951986e-10 luc = 8.885592091e-17 wuc = 2.592975112e-18 puc = -5.198338163e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.309699835e+05 lvsat = -1.018707309e+00 wvsat = -1.810156698e-02 pvsat = 3.628961420e-7   a0 = 1.975981626e+00 la0 = -1.026409245e-05 wa0 = -1.661863951e-07 pa0 = 3.331667456e-12   ags = 1.357626087e-01 lags = -4.505258039e-07 wags = -1.096312172e-08 pags = 2.197861975e-13   a1 = 0.0   a2 = 1.422460665e+00 la2 = -9.070829603e-06 wa2 = -1.611809675e-07 pa2 = 3.231319771e-12   b0 = 2.084009113e-07 lb0 = -3.628224494e-12 wb0 = -3.968180608e-14 pb0 = 7.955319199e-19   b1 = -6.567510453e-09 lb1 = 5.148289577e-14 wb1 = -1.128835647e-16 pb1 = 2.263064306e-21   keta = 6.859544784e-02 lketa = -9.068448402e-07 wketa = -1.635807123e-08 pketa = 3.279429314e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -3.154612309e-01 lpclm = 6.625012403e-06 wpclm = 1.171469302e-07 ppclm = -2.348535299e-12   pdiblc1 = 0.39   pdiblc2 = 7.397364563e-03 lpdiblc2 = -1.226965081e-07 wpdiblc2 = -2.612521092e-09 ppdiblc2 = 5.237523503e-14   pdiblcb = -0.225   drout = 0.56   pscbe1 = 5.213741541e+08 lpscbe1 = 5.585828268e+03 wpscbe1 = 1.326905439e+02 ppscbe1 = -2.660150168e-3   pscbe2 = 4.583062919e-09 lpscbe2 = 1.098129321e-13 wpscbe2 = 2.035453843e-15 ppscbe2 = -4.080632067e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -2.661533322e-10 lalpha0 = 5.335782120e-15 walpha0 = 9.481233384e-17 palpha0 = -1.900776336e-21   alpha1 = -2.661533322e-10 lalpha1 = 5.335782120e-15 walpha1 = 9.481233384e-17 palpha1 = -1.900776336e-21   beta0 = 1.018613997e+02 lbeta0 = -1.440661172e-03 wbeta0 = -2.559933014e-05 pbeta0 = 5.132096107e-10   agidl = 3.239573667e-09 lagidl = -2.685031118e-14 wagidl = -2.023356074e-16 pagidl = 4.056378731e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.976589972e-01 lkt1 = 3.195795709e-06 wkt1 = 7.298204048e-08 pkt1 = -1.463127527e-12   kt2 = -7.255181933e-02 lkt2 = 2.807855146e-07 wkt2 = 3.480389165e-09 pkt2 = -6.977405889e-14   at = -2.587278737e+04 lat = 1.941883367e+00 wat = 4.907651657e-02 pat = -9.838749621e-7   ute = 5.887236790e-01 lute = -1.346616422e-05 wute = -1.162380250e-08 pute = 2.330313772e-13   ua1 = 5.604456060e-09 lua1 = -7.045301479e-14 wua1 = -8.685606108e-16 pua1 = 1.741270770e-20   ub1 = -4.976686216e-18 lub1 = 7.513477481e-23 wub1 = 1.106512604e-24 pub1 = -2.218311572e-29   uc1 = -1.240647521e-10 luc1 = 1.890019067e-15 wuc1 = 1.401021188e-17 puc1 = -2.808735755e-22   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.182 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.225466592e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.268897418e-07 wvth0 = 4.029261970e-08 pvth0 = -3.580957367e-13   k1 = 5.173430238e-01 lk1 = 1.246276280e-08 wk1 = -2.709336663e-08 pk1 = -3.253459562e-14   k2 = -1.984361416e-02 lk2 = 2.435446056e-08 wk2 = 1.591907642e-08 pk2 = -1.128310244e-16   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-3.262144225e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.845186621e-07 wvoff = 4.036774869e-08 pvoff = -2.205396355e-13   nfactor = {2.749762786e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.230592494e-05 wnfactor = 3.428338356e-07 pnfactor = -3.632163080e-12   eta0 = 0.08   etab = -0.07   u0 = 2.569142681e-02 lu0 = -6.683398164e-08 wu0 = -7.707636664e-09 pu0 = 3.568482746e-14   ua = -2.645955641e-09 lua = 9.842667002e-15 wua = 7.959372975e-16 pua = -4.039427123e-21   ub = 7.945722027e-18 lub = -2.979053486e-23 wub = -3.082850868e-24 pub = 1.408506601e-29   uc = -9.000950918e-11 luc = -7.278918832e-17 wuc = -8.094321519e-18 puc = 3.402557702e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.225680401e+04 lvsat = 5.363384013e-01 wvsat = 5.986814741e-02 pvsat = -2.645865762e-7   a0 = 8.325157453e-02 la0 = 4.968173143e-06 wa0 = 5.170162854e-07 pa0 = -2.166593996e-12   ags = 5.468507736e-03 lags = 5.980518049e-07 wags = 1.851654966e-08 pags = -1.745956482e-14   a1 = 0.0   a2 = -2.153515568e-01 la2 = 4.109914648e-06 wa2 = 4.835429026e-07 pa2 = -1.957272872e-12   b0 = -2.605333648e-07 lb0 = 1.456530502e-13 wb0 = 8.213522359e-14 pb0 = -1.848241260e-19   b1 = 4.970262244e-09 lb1 = -4.137050290e-14 wb1 = -6.640762609e-16 pb1 = 6.698939107e-21   keta = -7.471031958e-02 lketa = 2.464477322e-07 wketa = 3.917160216e-08 pketa = -1.189473859e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -7.174366670e-01 lpclm = 9.860020268e-06 wpclm = 1.443821376e-07 ppclm = -2.567718120e-12   pdiblc1 = 0.39   pdiblc2 = -1.577993739e-02 lpdiblc2 = 6.382920311e-08 wpdiblc2 = 7.625047579e-09 ppdiblc2 = -3.001441418e-14   pdiblcb = -0.225   drout = 0.56   pscbe1 = 1.635877538e+09 lpscbe1 = -3.383444200e+03 wpscbe1 = -3.980716316e+02 ppscbe1 = 1.611304398e-3   pscbe2 = 2.885572840e-08 lpscbe2 = -8.552801828e-14 wpscbe2 = -6.764433676e-15 ppscbe2 = 3.001319411e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 7.984599966e-10 lalpha0 = -3.231986413e-15 walpha0 = -2.844370015e-16 palpha0 = 1.151336984e-21   alpha1 = 7.984599966e-10 lalpha1 = -3.231986413e-15 walpha1 = -2.844370015e-16 palpha1 = 1.151336984e-21   beta0 = -1.855841991e+02 lbeta0 = 8.726363315e-04 wbeta0 = 7.679799041e-05 pbeta0 = -3.108609856e-10   agidl = 2.708385822e-09 lagidl = -2.257543092e-14 wagidl = -9.585594279e-16 pagidl = 1.014229789e-20   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 1.241541157e-01 lkt1 = -2.613193816e-06 wkt1 = -2.561424417e-07 pkt1 = 1.185592253e-12   kt2 = -1.652854201e-02 lkt2 = -1.700772160e-07 wkt2 = -1.044116749e-08 pkt2 = 4.226349676e-14   at = 2.410983631e+05 lat = -2.066403835e-01 wat = -1.043107187e-01 pat = 2.505509955e-7   ute = -1.816653289e+00 lute = 5.891768405e-06 wute = -5.096625449e-08 pute = 5.496505787e-13   ua1 = -8.452568181e-09 lua1 = 4.267475348e-14 wua1 = 2.605681833e-15 pua1 = -1.054721378e-20   ub1 = 9.913264274e-18 lub1 = -4.469619649e-23 wub1 = -3.319537812e-24 pub1 = 1.343674217e-29   uc1 = 1.812655859e-09 luc1 = -1.369627265e-14 wuc1 = -5.976163336e-16 puc1 = 4.641359246e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.183 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-9.374971238e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.387458718e-07 wvth0 = -9.902393603e-08 pvth0 = 2.058263347e-13   k1 = 4.262586436e-01 lk1 = 3.811518396e-07 wk1 = -1.983617283e-08 pk1 = -6.191008326e-14   k2 = 5.828676888e-02 lk2 = -2.918997507e-07 wk2 = -7.619590015e-09 pk2 = 9.516639452e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.671662094e-01 ldsub = -1.243339703e-06 wdsub = 1.447513065e-14 pdsub = -5.859207253e-20   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-7.637682659e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.267677129e-07 wvoff = -6.652184573e-08 pvoff = 2.121253926e-13   nfactor = {3.460589021e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.887186817e-07 wnfactor = -5.926071800e-07 pnfactor = 1.542916771e-13   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411601813e-01 letab = 2.880404027e-7   u0 = -9.130858720e-04 lu0 = 4.085509968e-08 wu0 = 6.498323175e-09 pu0 = -2.181770163e-14   ua = 9.144852156e-10 lua = -4.569196486e-15 wua = -5.823619166e-16 pua = 1.539617978e-21   ub = -3.798981527e-18 lub = 1.774938256e-23 wub = 2.347864378e-24 pub = -7.897247394e-30   uc = -9.862164776e-11 luc = -3.792918907e-17 wuc = -1.690838641e-17 puc = 6.970292854e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.588091081e+05 lvsat = -3.584866709e-01 wvsat = -3.553530294e-02 pvsat = 1.215851250e-7   a0 = 1.735953108e+00 la0 = -1.721590805e-06 wa0 = -1.588941016e-07 pa0 = 5.693391711e-13   ags = -4.963517975e-01 lags = 2.629307491e-06 wags = 2.139736755e-07 pags = -8.086260323e-13   a1 = 0.0   a2 = 0.8   b0 = -2.798923892e-07 lb0 = 2.240140252e-13 wb0 = 3.996161075e-14 pb0 = -1.411483033e-20   b1 = 9.073726748e-08 lb1 = -3.885360425e-13 wb1 = -4.466338120e-14 pb1 = 1.847982257e-19   keta = 6.055649189e-03 lketa = -8.047473700e-08 wketa = 8.071242217e-09 pketa = 6.939873608e-15   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.269494961e+00 lpclm = -2.230406903e-06 wpclm = -7.926915954e-07 ppclm = 1.225345510e-12   pdiblc1 = 0.39   pdiblc2 = -5.085006988e-04 lpdiblc2 = 2.013863468e-09 wpdiblc2 = 4.414225528e-10 ppdiblc2 = -9.367163891e-16   pdiblcb = -1.037679986e+00 lpdiblcb = 3.289545732e-06 wpdiblcb = 2.895026170e-07 ppdiblcb = -1.171841455e-12   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 5.676192454e-09 lpscbe2 = 8.297527828e-15 wpscbe2 = 1.443812342e-15 ppscbe2 = -3.211938916e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.023887500e-10 lalpha0 = 4.144466225e-16   alpha1 = -1.023887500e-10 lalpha1 = 4.144466225e-16   beta0 = 5.212771198e+01 lbeta0 = -8.956799935e-05 wbeta0 = 1.375364980e-06 pbeta0 = -5.567167980e-12   agidl = -3.216199767e-09 lagidl = 1.405958515e-15 wagidl = 1.494070646e-15 pagidl = 2.146031928e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -8.444312620e-01 lkt1 = 1.307421861e-06 wkt1 = 1.947823037e-07 pkt1 = -6.396496584e-13   kt2 = -5.808477657e-02 lkt2 = -1.866928689e-09 wkt2 = -2.468009810e-09 pkt2 = 9.989948407e-15   at = 2.523242358e+05 lat = -2.520801905e-01 wat = -4.235147391e-02 pat = -2.460867056e-10   ute = -2.859903611e+00 lute = 1.011461098e-05 wute = 1.318901819e-06 pute = -4.995267164e-12   ua1 = 3.219835857e-10 lua1 = 7.157342196e-15 wua1 = 1.226072533e-15 pua1 = -4.962865747e-21   ub1 = -1.641079922e-18 lub1 = 2.073189084e-24 wub1 = -1.300301004e-25 pub1 = 5.263325897e-31   uc1 = -3.165394879e-09 luc1 = 6.453756676e-15 wuc1 = 1.087119518e-15 puc1 = -2.178072417e-21   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.184 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.064238990e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.792070468e-07 wvth0 = -4.382037523e-08 pvth0 = 9.278186294e-14   k1 = 6.368438488e-01 lk1 = -5.007927892e-08 wk1 = -6.209934803e-08 pk1 = 2.463539035e-14   k2 = -5.155586817e-02 lk2 = -6.696674458e-08 wk2 = 2.332659811e-08 pk2 = 3.179556413e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 2.561714481e+00 ldsub = -4.713393291e-06 wdsub = -1.096150081e-06 pdsub = 2.244668703e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.659232465e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.433967928e-07 wvoff = -2.075543970e-08 pvoff = 1.184060905e-13   nfactor = {2.779446446e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.061080548e-07 wnfactor = -1.294881637e-07 pnfactor = -7.940718665e-13   eta0 = -1.352200576e+00 leta0 = 2.770026422e-06 weta0 = 3.999466407e-07 peta0 = -8.190007321e-13   etab = -2.628395144e+00 letab = 5.381337978e-06 wetab = 1.251860488e-06 petab = -2.563528610e-12   u0 = 2.538673143e-02 lu0 = -1.300100868e-08 wu0 = -5.902161450e-09 pu0 = 3.575700776e-15   ua = 5.420902728e-10 lua = -3.806615432e-15 wua = -4.410015722e-16 pua = 1.250143799e-21   ub = 3.919589790e-18 lub = 1.943485184e-24 wub = -1.174438393e-24 pub = -6.843638367e-31   uc = -2.265406637e-10 luc = 2.240201737e-16 wuc = 5.047201046e-17 puc = -6.827696366e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.235242104e+05 lvsat = 2.196684404e-01 wvsat = 6.593974298e-02 pvsat = -8.621293713e-8   a0 = 1.189678917e-01 la0 = 1.589631096e-06 wa0 = 4.330178381e-07 pa0 = -6.427633012e-13   ags = 1.764897963e+00 lags = -2.001223237e-06 wags = -7.244085993e-07 pags = 1.112969731e-12   a1 = 0.0   a2 = 0.8   b0 = 3.906020074e-07 lb0 = -1.149007638e-12 wb0 = -1.892066835e-13 pb0 = 4.551702735e-19   b1 = -2.192794395e-07 lb1 = 2.463084197e-13 wb1 = 1.011754364e-13 pb1 = -1.138468590e-19   keta = -1.069478165e-01 lketa = 1.509309349e-07 wketa = 4.249823647e-08 pketa = -6.355886455e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.055608415e+00 lpclm = 2.553596197e-07 wpclm = -6.295432144e-08 ppclm = -2.689922364e-13   pdiblc1 = 4.093380786e-01 lpdiblc1 = -3.960003384e-08 wpdiblc1 = -6.384733359e-09 ppdiblc1 = 1.307449735e-14   pdiblc2 = 5.220251998e-04 lpdiblc2 = -9.642170375e-11 wpdiblc2 = -3.278232098e-11 ppdiblc2 = 3.434849637e-17   pdiblcb = 1.400359973e+00 lpdiblcb = -1.703011546e-06 wpdiblcb = -5.790052339e-07 ppdiblcb = 6.066672090e-13   drout = 7.123697981e-01 ldrout = -3.120190633e-07 wdrout = -1.605669185e-07 pdrout = 3.288049216e-13   pscbe1 = 800000000.0   pscbe2 = 1.008053695e-08 lpscbe2 = -7.215787272e-16 wpscbe2 = -1.446915996e-16 ppscbe2 = 4.095974328e-23   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.813025868e-11 lalpha0 = 1.471730595e-16 walpha0 = 3.422667065e-17 palpha0 = -7.008852048e-23   alpha1 = -5.220849730e-10 lalpha1 = 1.273890056e-15 walpha1 = 2.962567709e-16 palpha1 = -6.066672090e-22   beta0 = 9.742426847e+00 lbeta0 = -2.772472095e-06 wbeta0 = -2.438830683e-06 pbeta0 = 2.243446542e-12   agidl = -6.909725199e-09 lagidl = 8.969467556e-15 wagidl = 3.482029897e-15 pagidl = -3.856290063e-21   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 1.300435457e-01 lkt1 = -6.880832881e-07 wkt1 = -2.645313280e-07 pkt1 = 3.009213137e-13   kt2 = -7.872188383e-02 lkt2 = 4.039322364e-08 wkt2 = 9.121859679e-09 pkt2 = -1.374349658e-14   at = 1.730672227e+05 lat = -8.977966041e-02 wat = -6.919883191e-02 pat = 5.473126182e-8   ute = 5.476344856e+00 lute = -6.956150226e-06 wute = -2.351571000e-06 pute = 2.521035313e-12   ua1 = 7.715539567e-09 lua1 = -7.982996903e-15 wua1 = -2.189208279e-15 pua1 = 2.030860918e-21   ub1 = -1.238420084e-18 lub1 = 1.248632333e-24 wub1 = -1.898271103e-25 pub1 = 6.487834116e-31   uc1 = 2.666721875e-11 luc1 = -8.286828639e-17 wuc1 = -1.144566031e-17 puc1 = 7.154189188e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.185 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.353572138e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.239489920e-07 wvth0 = 7.794876132e-08 pvth0 = -3.480479412e-14   k1 = 9.698768557e-01 lk1 = -3.990229377e-07 wk1 = -1.818242934e-07 pk1 = 1.500801949e-13   k2 = -2.801694580e-01 lk2 = 1.725688595e-07 wk2 = 1.115937703e-07 pk2 = -6.068857217e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -7.560800600e+00 ldsub = 5.892724949e-06 wdsub = 3.338430896e-06 pdsub = -2.401774379e-12   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-5.367594122e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.451560707e-07 wvoff = 1.364086522e-07 pvoff = -4.626651584e-14   nfactor = {8.348410593e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.028913354e-06 wnfactor = -2.850370582e-06 pnfactor = 2.056800709e-12   eta0 = 4.264527448e+00 leta0 = -3.115040783e-06 weta0 = -1.546162993e-06 peta0 = 1.220084289e-12   etab = 5.259069981e+00 letab = -2.882950793e-06 wetab = -2.505260119e-06 petab = 1.373088434e-12   u0 = 1.115496045e-02 lu0 = 1.910685152e-09 wu0 = -1.089516501e-09 pu0 = -1.466868285e-15   ua = -9.014773405e-09 lua = 6.206827408e-15 wua = 3.036833109e-15 pua = -2.393844434e-21   ub = 1.456060757e-17 lub = -9.205907223e-24 wub = -5.055593347e-24 pub = 3.382213296e-30   uc = 1.264062873e-10 luc = -1.457888178e-16 wuc = -7.847839194e-17 puc = 6.683404421e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -2.863805546e+04 lvsat = 1.202490994e-01 wvsat = 1.148198481e-02 pvsat = -2.915345957e-8   a0 = 1.323171951e+00 la0 = 3.278961875e-07 wa0 = 4.316925212e-08 pa0 = -2.342896990e-13   ags = -1.673452048e+00 lags = 1.601393945e-06 wags = 7.079050207e-07 pags = -3.877726727e-13   a1 = 0.0   a2 = 2.691326384e+00 la2 = -1.981684502e-06 wa2 = -7.400968748e-07 pa2 = 7.754550030e-13   b0 = -1.479489239e-06 lb0 = 8.104272180e-13 wb0 = 5.138484814e-13 pb0 = -2.814733519e-19   b1 = 3.310580984e-08 lb1 = -1.813453499e-14 wb1 = -1.567553233e-14 pb1 = 8.586664725e-21   keta = 1.721419199e-01 lketa = -1.414923137e-07 wketa = -6.030256514e-08 pketa = 4.415324536e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 9.689395440e-01 lpclm = 3.461690957e-07 wpclm = -6.031833415e-08 ppclm = -2.717541580e-13   pdiblc1 = 5.171917665e-01 lpdiblc1 = -1.526064317e-07 wpdiblc1 = 1.007999859e-07 ppdiblc1 = -9.923097187e-14   pdiblc2 = -2.505533020e-03 lpdiblc2 = 3.075778110e-09 wpdiblc2 = 1.203058380e-09 ppdiblc2 = -1.260534494e-15   pdiblcb = 1.812254072e-01 lpdiblcb = -4.256328260e-07 wpdiblcb = -1.934575381e-07 ppdiblcb = 2.026999720e-13   drout = 1.895053150e+00 ldrout = -1.551205112e-06 wdrout = -4.347315981e-07 pdrout = 6.160678188e-13   pscbe1 = 3.677005472e+09 lpscbe1 = -3.014454409e+03 wpscbe1 = -1.024881413e+03 ppscbe1 = 1.073845123e-3   pscbe2 = -2.904556904e-07 lpscbe2 = 3.141727669e-13 wpscbe2 = 1.066891464e-13 ppscbe2 = -1.118968649e-19   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 2.437394826e-10 lalpha0 = -7.873689510e-17 walpha0 = -6.845334129e-17 palpha0 = 3.749702903e-23   alpha1 = 1.344169946e-09 lalpha1 = -6.815251922e-16 walpha1 = -5.925135417e-16 palpha1 = 3.245641053e-22   beta0 = 4.724384272e+00 lbeta0 = 2.485307465e-06 wbeta0 = -1.963094245e-07 pbeta0 = -1.062111692e-13   agidl = 2.739012397e-09 lagidl = -1.140238478e-15 wagidl = -5.493592103e-16 pagidl = 3.676986587e-22   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -6.385840845e-01 lkt1 = 1.172655272e-07 wkt1 = 7.848051081e-08 pkt1 = -5.847791574e-14   kt2 = -1.894576718e-02 lkt2 = -2.223869698e-08 wkt2 = -8.371680120e-09 pkt2 = 4.585797078e-15   at = 9.546769770e+04 lat = -8.472818105e-03 wat = -3.554708856e-02 pat = 1.947180643e-8   ute = -1.947290279e+00 lute = 8.221490771e-07 wute = 5.818240792e-09 pute = 5.102180192e-14   ua1 = -2.740241179e-09 lua1 = 2.972308768e-15 wua1 = 6.457714406e-18 pua1 = -2.697030184e-22   ub1 = 1.073873251e-18 lub1 = -1.174130816e-24 wub1 = 7.937885005e-25 pub1 = -3.818244350e-31   uc1 = -3.606988557e-11 luc1 = -1.713391691e-17 wuc1 = 1.190988303e-16 puc1 = -6.523936176e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.186 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.085259194e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.302613092e-08 wvth0 = -1.768630066e-08 pvth0 = 1.758170196e-14   k1 = 8.087701363e-01 lk1 = -3.107727045e-07 wk1 = -2.590948188e-07 pk1 = 1.924070570e-13   k2 = -2.145098705e-01 lk2 = 1.366021790e-07 wk2 = 1.589852737e-07 pk2 = -8.664845295e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 5.636914301e+00 ldsub = -1.336653331e-06 wdsub = -2.086058300e-06 pdsub = 5.696251895e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.681786805e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.674323964e-08 wvoff = 2.443840692e-08 pvoff = 1.506798525e-14   nfactor = {-6.089441816e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.879781249e-06 wnfactor = 2.742384338e-06 pnfactor = -1.006770617e-12   eta0 = -3.699796044e+00 leta0 = 1.247616518e-06 weta0 = 1.492539424e-06 peta0 = -4.444409273e-13   etab = -8.337616450e-03 letab = 2.403403592e-09 wetab = 2.967899333e-09 petab = -8.561692685e-16   u0 = 1.278396954e-02 lu0 = 1.018354697e-09 wu0 = -2.008454712e-09 pu0 = -9.634969070e-16   ua = -5.382351371e-10 lua = 1.563591658e-15 wua = 2.360190453e-16 pua = -8.596285104e-22   ub = 4.927081914e-19 lub = -1.499863640e-24 wub = -4.515736510e-25 pub = 8.602464067e-31   uc = -3.005952652e-10 luc = 8.811195762e-17 wuc = 9.328092264e-17 puc = -2.725141434e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.379014284e+05 lvsat = -8.053206641e-02 wvsat = -1.261133885e-01 pvsat = 4.621784607e-8   a0 = 5.428872036e+00 la0 = -1.921103676e-06 wa0 = -1.771368292e-06 pa0 = 7.596686045e-13   ags = 3.777282979e-02 lags = 6.640277382e-07 wags = 4.318341093e-07 pags = -2.365479292e-13   a1 = 0.0   a2 = -4.192587869e+00 la2 = 1.789151628e-06 wa2 = 2.058660077e-06 pa2 = -7.576340860e-13   b0 = 0.0   b1 = 0.0   keta = -1.385779520e-01 lketa = 2.871226418e-08 wketa = 3.857065034e-08 pketa = -1.000703025e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 3.418654332e+00 lpclm = -9.957234223e-07 wpclm = -1.538210267e-06 ppclm = 5.377980956e-13   pdiblc1 = -7.259627459e-01 lpdiblc1 = 5.283625313e-07 wpdiblc1 = 1.891142993e-07 ppdiblc1 = -1.476073449e-13   pdiblc2 = -1.005717226e-02 lpdiblc2 = 7.212377295e-09 wpdiblc2 = 7.631729514e-10 ppdiblc2 = -1.019576253e-15   pdiblcb = -7.395560085e-01 lpdiblcb = 7.874821395e-08 wpdiblcb = 2.807954137e-07 ppdiblcb = -5.708393870e-14   drout = -1.022448742e+00 ldrout = 4.692948698e-08 wdrout = 7.212653210e-07 pdrout = -1.715839361e-14   pscbe1 = -4.953995917e+09 lpscbe1 = 1.713392377e+03 wpscbe1 = 2.049770818e+03 ppscbe1 = -6.103725031e-4   pscbe2 = 6.114103046e-07 lpscbe2 = -1.798468785e-13 wpscbe2 = -2.146169615e-13 ppscbe2 = 6.410658839e-20   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.029992194e+01 lbeta0 = -5.688326813e-07 wbeta0 = -1.150113866e-06 pbeta0 = 4.162590589e-13   agidl = 1.179342156e-08 lagidl = -6.100017458e-15 wagidl = -4.662590850e-15 pagidl = 2.620824120e-21   bgidl = -1.369778406e+08 lbgidl = 6.228080366e+02 wbgidl = 4.050278901e+02 pbgidl = -2.218641525e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.727537085e-01 lkt1 = -2.834970704e-08 wkt1 = -3.091015358e-08 pkt1 = 1.443555441e-15   kt2 = -3.050418753e-02 lkt2 = -1.590728327e-08 wkt2 = -1.764767435e-08 pkt2 = 9.666954815e-15   at = 2.257973119e+05 lat = -7.986412251e-02 wat = -6.256276301e-02 pat = 3.427031751e-8   ute = 1.464124599e+00 lute = -1.046538708e-06 wute = -4.728234654e-07 pute = 3.132097625e-13   ua1 = 5.527642041e-09 lua1 = -1.556630963e-15 wua1 = -1.061789486e-15 pua1 = 3.154560918e-22   ub1 = -1.350208997e-18 lub1 = 1.537208377e-25 wub1 = -1.650472036e-25 pub1 = 1.434017928e-31   uc1 = 1.088720582e-10 luc1 = -9.652949014e-17 wuc1 = -6.660029172e-17 puc1 = 3.648197480e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.187 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.173288692e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.186853037e-09 wvth0 = 4.516975170e-08 pvth0 = -1.135259031e-15   k1 = -6.612031822e+00 lk1 = 1.898956599e-06 wk1 = 2.658800115e-06 pk1 = -6.764691070e-13   k2 = 2.514527904e+00 lk2 = -6.760370444e-07 wk2 = -9.407527209e-07 pk2 = 2.408260284e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 5.675709544e+00 ldsub = -1.348205585e-06 wdsub = -1.785995441e-06 pdsub = 4.802739718e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.154781360e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.265864425e-08 wvoff = 2.400724609e-08 pvoff = 1.519637416e-14   nfactor = {1.349410693e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.951709977e-06 wnfactor = -4.169761294e-06 pnfactor = 1.051493549e-12   eta0 = 4.900000033e-01 leta0 = -3.431226414e-16 weta0 = -1.166378993e-15 peta0 = 1.222312251e-22   etab = 9.805127857e-03 letab = -2.999052094e-09 wetab = -3.495126757e-09 petab = 1.068358325e-15   u0 = 5.003295632e-02 lu0 = -1.007346234e-08 wu0 = -1.729511929e-08 pu0 = 3.588489637e-15   ua = 2.206544280e-08 lua = -5.167218539e-15 wua = -8.832428961e-15 pua = 1.840728595e-21   ub = -1.961024278e-17 lub = 4.486292587e-24 wub = 7.804349067e-24 pub = -1.598160981e-30   uc = 1.546925540e-10 luc = -4.746137276e-17 wuc = -5.501451545e-17 puc = 1.690725974e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 8.065087060e+05 lvsat = -2.200715985e-01 wvsat = -2.341771938e-01 pvsat = 7.839654568e-8   a0 = -4.411010424e+00 la0 = 1.008967323e-06 wa0 = 1.986821790e-06 pa0 = -3.594264474e-13   ags = 5.579382640e+00 lags = -9.861251231e-07 wags = -1.542264637e-06 pags = 3.512893249e-13   a1 = 0.0   a2 = 2.426986337e+00 la2 = -1.819920811e-07 wa2 = -7.033766595e-07 pa2 = 6.483140305e-14   b0 = 0.0   b1 = 0.0   keta = -2.897652166e-01 lketa = 7.373205188e-08 wketa = 9.317122479e-08 pketa = -2.626571631e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.869351875e-01 lpclm = -6.317575404e-08 wpclm = 1.922670072e-07 ppclm = 2.250522521e-14   pdiblc1 = 1.688364233e+00 lpdiblc1 = -1.905636848e-07 wpdiblc1 = -5.345603795e-07 ppdiblc1 = 6.788488258e-14   pdiblc2 = 1.089412085e-01 lpdiblc2 = -2.822236553e-08 wpdiblc2 = -3.642358206e-08 ppdiblc2 = 1.005370972e-14   pdiblcb = 1.051487354e+01 lpdiblcb = -3.272539544e-06 wpdiblcb = -3.825886630e-06 ppdiblcb = 1.165783307e-12   drout = -6.951243309e+00 ldrout = 1.812376289e-06 wdrout = 2.831811997e-06 pdrout = -6.456264302e-13   pscbe1 = 7.996425337e+08 lpscbe1 = 1.026875649e-01 wpscbe1 = 1.161374235e-01 ppscbe1 = -3.658059663e-8   pscbe2 = 5.509424902e-08 lpscbe2 = -1.418986507e-14 wpscbe2 = -1.630714916e-14 ppscbe2 = 5.054884015e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 1.556957958e+01 lbeta0 = -2.138004986e-06 wbeta0 = -2.309938342e-06 pbeta0 = 7.616257922e-13   agidl = -2.207792597e-08 lagidl = 3.986023054e-15 wagidl = 8.907296094e-15 pagidl = -1.419948965e-21   bgidl = 5.060634582e+09 lbgidl = -9.249110024e+02 wbgidl = -1.446527978e+03 pbgidl = 3.294828962e-4   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 3.585729792e-01 lkt1 = -2.461205115e-07 wkt1 = -3.204994294e-07 pkt1 = 8.767600204e-14   kt2 = -1.101023874e-01 lkt2 = 7.795070678e-09 wkt2 = 2.414162440e-08 pkt2 = -2.776853618e-15   at = 5.982053422e+05 lat = -1.907579237e-01 wat = -1.756809199e-01 pat = 6.795407669e-8   ute = -6.587427353e+00 lute = 1.351012175e-06 wute = 2.195243134e-06 pute = -4.812737691e-13   ua1 = -4.094201923e-10 lua1 = 2.112777436e-16 wua1 = 2.503421065e-16 pua1 = -7.526389315e-23   ub1 = -1.550050639e-18 lub1 = 2.132286827e-25 wub1 = 5.716186444e-25 pub1 = -7.595888011e-32   uc1 = -1.100972588e-09 luc1 = 2.637319995e-16 wuc1 = 3.714208734e-16 puc1 = -9.394977764e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.188 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.4e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.533757844e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.165854072e-08 wvth0 = 2.877864694e-07 pvth0 = -6.060649623e-14   k1 = 5.024837192e+00 lk1 = -8.077292811e-07 wk1 = -1.793602667e-06 pk1 = 3.628794740e-13   k2 = -1.203945379e+00 lk2 = 1.836961905e-07 wk2 = 5.683154989e-07 pk2 = -1.105820809e-13   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -7.140496224e-02 ldsub = -4.207903137e-08 wdsub = 7.082498285e-07 pdsub = -9.440963904e-14   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {1.114141508e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.713001229e-07 wvoff = -3.467769597e-07 pvoff = 1.070892604e-13   nfactor = {-2.314243600e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.795698776e-06 wnfactor = 8.641330019e-06 pnfactor = -2.005863047e-12   eta0 = 8.637332848e+00 leta0 = -1.994263397e-06 weta0 = -2.902340675e-06 peta0 = 7.104204386e-13   etab = 4.457350556e-01 letab = -1.099276346e-07 wetab = -1.572093036e-07 petab = 3.877348296e-14   u0 = 2.772128615e-02 lu0 = -5.363956707e-09 wu0 = -1.287528550e-08 pu0 = 2.774451949e-15   ua = 1.559585230e-08 lua = -3.969280173e-15 wua = -8.521885237e-15 pua = 1.902098137e-21   ub = -2.444535102e-17 lub = 6.004640905e-24 wub = 1.164490698e-23 pub = -2.657512380e-30   uc = -8.134594543e-10 luc = 1.859757529e-16 wuc = 3.393974039e-16 puc = -7.837304353e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -6.166334752e+06 lvsat = 1.470281103e+00 wvsat = 2.370845596e+00 pvsat = -5.533967770e-7   a0 = -7.262363205e+00 la0 = 1.782211533e-06 wa0 = 3.414027580e-06 pa0 = -7.355965577e-13   ags = 1.250000289e+00 lags = -6.250419382e-14 wags = -1.030797581e-13 pags = 2.226599349e-20   a1 = 0.0   a2 = 1.204164765e-01 la2 = 3.690155671e-07 wa2 = -3.449132912e-07 pa2 = -1.807277248e-14   b0 = 2.304770800e-06 lb0 = -5.641502725e-13 wb0 = -8.210331115e-13 pb0 = 2.009683799e-19   b1 = 0.0   keta = -1.157229628e+00 lketa = 2.915686491e-07 wketa = 3.741828346e-07 pketa = -9.701067631e-14   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -4.322075013e+00 lpclm = 1.060279592e-06 wpclm = 2.349533807e-06 ppclm = -5.038600769e-13   pdiblc1 = 5.546902471e+00 lpdiblc1 = -1.149260113e-06 wpdiblc1 = -1.846554770e-06 ppdiblc1 = 3.940949015e-13   pdiblc2 = -1.061694132e-01 lpdiblc2 = 2.232495904e-08 wpdiblc2 = 4.782757595e-08 ppdiblc2 = -9.818508289e-15   pdiblcb = -3.933633725e+01 lpdiblcb = 8.685544401e-06 wpdiblcb = 1.464998859e-05 ppdiblcb = -3.269640747e-12   drout = 1.045917173e+00 ldrout = -9.861861236e-09 wdrout = -2.186712514e-08 pdrout = 4.696511932e-15   pscbe1 = 1.315112124e+09 lpscbe1 = -1.260637174e+02 wpscbe1 = -1.835897369e+02 ppscbe1 = 4.492729458e-5   pscbe2 = -1.189011271e-07 lpscbe2 = 2.734079173e-14 wpscbe2 = 4.528227468e-14 ppscbe2 = -9.643395651e-21   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 8.537401523e-01 lbeta0 = 1.304494488e-06 wbeta0 = 4.725869381e-06 pbeta0 = -9.037200591e-13   agidl = 5.062513637e-08 lagidl = -1.351237198e-14 wagidl = -2.008634739e-14 pagidl = 5.570992149e-21   bgidl = 1.000001405e+09 lbgidl = -3.014149466e-04 wbgidl = -5.003471642e-04 pbgidl = 1.073736496e-10   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -8.137015679e-01 lkt1 = 2.245377252e-08 wkt1 = 4.869712264e-08 pkt1 = 3.849619390e-15   kt2 = 9.165548643e-01 lkt2 = -2.429231726e-07 wkt2 = -3.251522521e-07 pkt2 = 8.251430439e-14   at = -2.715579333e+06 lat = 6.061364917e-01 wat = 1.177939287e+00 pat = -2.583065531e-7   ute = -4.184706860e+00 lute = 8.637191361e-07 wute = 6.715658060e-07 pute = -1.442355461e-13   ua1 = 8.654142657e-10 lua1 = -8.500113454e-17 wua1 = -1.607646214e-15 pua1 = 3.739078732e-22   ub1 = -2.367243183e-20 lub1 = -1.444762082e-25 wub1 = 1.772458897e-24 pub1 = -3.755637484e-31   uc1 = -4.959628665e-11 luc1 = 2.606501791e-17 wuc1 = 5.925262012e-17 puc1 = -2.455074041e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.189 pmos  lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.132197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.43165561   k2 = 0.041298226   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 3.2465718e-7   voff = {-0.18331232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7163132+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.08   etab = -0.07   u0 = 0.00786119   ua = -7.1939916e-10   ub = 6.0823395e-19   uc = -1.0566299e-10   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.464   ags = 0.11329   a1 = 0.0   a2 = 0.97   b0 = 2.7422e-8   b1 = -3.9995e-9   keta = 0.023361259   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.015   pdiblc1 = 0.39   pdiblc2 = 0.0012771588   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 1.0060625e-8   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.9002574e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.43825   kt2 = -0.058546   at = 70990.0   ute = -0.08298   ua1 = 2.0902e-9   ub1 = -1.2289e-18   uc1 = -2.9789e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.190 pmos  lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.122306285e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.982868384e-7   k1 = 4.317681715e-01 lk1 = -2.256608555e-9   k2 = 5.033022846e-02 lk2 = -1.810715531e-7   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = -6.164091325e-06 lcit = 1.300849701e-10 wcit = -2.117582368e-28 pcit = -8.470329473e-33   voff = {-1.605913386e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.555051222e-7   nfactor = {1.861696457e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.914610816e-6   eta0 = 0.08   etab = -0.07   u0 = 7.635644399e-03 lu0 = 4.521687458e-9   ua = -8.010813065e-10 lua = 1.637545294e-15   ub = 6.788117698e-19 lub = -1.414928252e-24   uc = -1.028163042e-10 luc = -5.706971639e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 80156.0   a0 = 1.509469929e+00 la0 = -9.115709008e-7   ags = 1.049873788e-01 lags = 1.664490819e-7   a1 = 0.0   a2 = 0.97   b0 = 9.700775719e-08 lb0 = -1.395039603e-12 wb0 = 1.323488980e-29   b1 = -6.884392611e-09 lb1 = 5.783567796e-14   keta = 2.267573477e-02 lketa = 1.374323550e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 1.338887300e-02 lpclm = 3.229951157e-8   pdiblc1 = 0.39   pdiblc2 = 6.360147655e-05 lpdiblc2 = 2.432912417e-8   pdiblcb = -0.225   drout = 0.56   pscbe1 = 8.938576588e+08 lpscbe1 = -1.881637226e+3   pscbe2 = 1.029690627e-08 lpscbe2 = -4.736913650e-15 wpscbe2 = 3.308722450e-30   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 2.671585369e-09 lagidl = -1.546340958e-14   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -3.927867777e-01 lkt1 = -9.114364509e-7   kt2 = -6.278181224e-02 lkt2 = 8.491861076e-8   at = 1.118928164e+05 lat = -8.200104608e-1   ute = 5.560938128e-01 lute = -1.281200801e-05 pute = 6.661338148e-28   ua1 = 3.166267995e-09 lua1 = -2.157276905e-14   ub1 = -1.870528981e-18 lub1 = 1.286323345e-23   uc1 = -8.473585446e-11 luc1 = 1.101562175e-15 wuc1 = 1.292469707e-32 puc1 = 2.067951531e-37   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.191 pmos  lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.112358787e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.783420642e-7   k1 = 4.412876255e-01 lk1 = -7.886703245e-8   k2 = 2.484377053e-02 lk2 = 2.403772589e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.56   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.128957182e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.457124407e-8   nfactor = {1.237365496e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.109864282e-6   eta0 = 0.08   etab = -0.07   u0 = 4.054862256e-03 lu0 = 3.333901647e-8   ua = -4.116327910e-10 lua = -1.496648732e-15   ub = -7.083317014e-19 lub = 9.748490297e-24 pub = -1.540743956e-45   uc = -1.127315598e-10 luc = 2.272602934e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 1.058026275e+05 lvsat = -2.063982878e-1   a0 = 1.534598689e+00 la0 = -1.113801512e-6   ags = 5.744741379e-02 lags = 5.490400238e-7   a1 = 0.0   a2 = 1.142030438e+00 la2 = -1.384462254e-6   b0 = -2.996670154e-08 lb0 = -3.731777287e-13   b1 = 3.106094340e-09 lb1 = -2.256551316e-14 wb1 = 2.067951531e-31 pb1 = 3.308722450e-36   keta = 3.525061082e-02 lketa = -8.745653760e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -3.121329953e-01 lpclm = 2.652026265e-06 ppclm = 1.942890293e-28   pdiblc1 = 0.39   pdiblc2 = 5.624786443e-03 lpdiblc2 = -2.042604117e-8   pdiblcb = -0.225   drout = 0.56   pscbe1 = 5.184270236e+08 lpscbe1 = 1.139744055e+3   pscbe2 = 9.866884960e-09 lpscbe2 = -1.276198935e-15   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 0.0   alpha1 = 0.0   beta0 = 30.0   agidl = 1.755673318e-11 lagidl = 5.895615726e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -5.948785418e-01 lkt1 = 7.149525958e-07 wkt1 = 2.220446049e-22   kt2 = -4.583856328e-02 lkt2 = -5.143684469e-8   at = -5.171844931e+04 lat = 4.966961934e-01 wat = 7.275957614e-18 pat = 2.910383046e-23   ute = -1.959723688e+00 lute = 7.434725183e-6   ua1 = -1.138003986e-09 lua1 = 1.306704339e-14 pua1 = -8.271806126e-37   ub1 = 5.947925689e-19 lub1 = -6.977119688e-24   uc1 = 1.350515634e-10 luc1 = -6.672375114e-16 wuc1 = 2.584939414e-32   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.192 pmos  lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.215473095e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.390414541e-7   k1 = 3.705753450e-01 lk1 = 2.073603688e-7   k2 = 3.689736530e-02 lk2 = -2.475251370e-08 wk2 = 1.387778781e-23   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 8.671662500e-01 ldsub = -1.243339868e-6   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.631142498e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.687020726e-7   nfactor = {1.797046218e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.555973533e-7   eta0 = 1.613990563e-01 leta0 = -3.294850649e-7   etab = -1.411601813e-01 letab = 2.880404027e-7   u0 = 1.732874298e-02 lu0 = -2.039066607e-8   ua = -7.202975006e-10 lua = -2.472434376e-16   ub = 2.791847984e-18 lub = -4.419449529e-24   uc = -1.460861833e-10 luc = 1.577380405e-16   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 5.905584912e+04 lvsat = -1.717784684e-2   a0 = 1.289912040e+00 la0 = -1.233650106e-7   ags = 1.043064125e-01 lags = 3.593653402e-7   a1 = 0.0   a2 = 0.8   b0 = -1.677137788e-07 lb0 = 1.843914468e-13 wb0 = 5.293955920e-29   b1 = -3.463996197e-08 lb1 = 1.302220299e-13 wb1 = 6.617444900e-30 pb1 = 3.308722450e-36   keta = 2.871291248e-02 lketa = -6.099340571e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 4.428331434e-02 lpclm = 1.209333237e-6   pdiblc1 = 0.39   pdiblc2 = 7.306427605e-04 lpdiblc2 = -6.156487289e-10   pdiblcb = -0.225   drout = 0.56   pscbe1 = 800000000.0   pscbe2 = 9.729203811e-09 lpscbe2 = -7.188966248e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = -1.023887500e-10 lalpha0 = 4.144466225e-16   alpha1 = -1.023887500e-10 lalpha1 = 4.144466225e-16   beta0 = 5.598858068e+01 lbeta0 = -1.051959272e-4   agidl = 9.778946584e-10 lagidl = 2.008383880e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -2.976462914e-01 lkt1 = -4.881766767e-7   kt2 = -6.501287345e-02 lkt2 = 2.617644868e-8   at = 1.334368986e+05 lat = -2.527709951e-1   ute = 8.424640015e-01 lute = -3.907900093e-06 wute = 1.110223025e-22 pute = -4.440892099e-28   ua1 = 3.763764597e-09 lua1 = -6.774212935e-15   ub1 = -2.006095138e-18 lub1 = 3.550688549e-24   uc1 = -1.136771268e-10 luc1 = 3.395602623e-16 wuc1 = -1.292469707e-32 puc1 = 2.584939414e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 3.0e-6   sbref = 3.0e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.193 pmos  lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.187249767e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.124642997e-8   k1 = 4.625210816e-01 lk1 = 1.907618818e-8   k2 = 1.392561050e-02 lk2 = 2.228847150e-8   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -5.153535000e-01 ldsub = 1.587749513e-06 pdsub = -1.110223025e-28   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.241870738e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.898797475e-8   nfactor = {2.415952533e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.422978233e-6   eta0 = -2.294866125e-01 leta0 = 4.709608354e-07 weta0 = 1.344410694e-23 peta0 = -1.994931997e-29   etab = 8.857767662e-01 letab = -1.814895405e-06 wetab = -1.344410694e-23 petab = 1.309716224e-28   u0 = 8.818423554e-03 lu0 = -2.963446712e-9   ua = -6.958714270e-10 lua = -2.972625406e-16   ub = 6.227540409e-19 lub = 2.236682050e-26   uc = -8.485768610e-11 luc = 3.235585476e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 6.157915752e+04 lvsat = -2.234501469e-2   a0 = 1.334517977e+00 la0 = -2.147079337e-7   ags = -2.686324314e-01 lags = 1.123060181e-6   a1 = 0.0   a2 = 0.8   b0 = -1.405313089e-07 lb0 = 1.287278646e-13   b1 = 6.473613569e-08 lb1 = -7.327785846e-14   keta = 1.235150666e-02 lketa = -2.748892790e-08 wketa = -8.673617380e-25 pketa = 8.673617380e-31   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 8.788856008e-01 lpclm = -4.997444597e-7   pdiblc1 = 3.914151144e-01 lpdiblc1 = -2.897835967e-9   pdiblc2 = 0.00043   pdiblcb = -0.225   drout = 2.616328668e-01 ldrout = 6.109887562e-7   pscbe1 = 800000000.0   pscbe2 = 9.674364571e-09 lpscbe2 = -6.065981997e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.242099782e-10 lalpha0 = -4.957658813e-17   alpha1 = 3.095550000e-10 lalpha1 = -4.291214901e-16 walpha1 = 5.169878828e-32   beta0 = 2.896240422e+00 lbeta0 = 3.525239907e-6   agidl = 2.864887684e-09 lagidl = -1.855753263e-15 wagidl = -8.271806126e-31   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -6.125380528e-01 lkt1 = 1.566508000e-7   kt2 = -5.311536987e-02 lkt2 = 1.813038296e-9   at = -2.118492732e+04 lat = 6.385971455e-02 pat = 7.275957614e-24   ute = -1.124889732e+00 lute = 1.207976995e-7   ua1 = 1.570083012e-09 lua1 = -2.282046628e-15 pua1 = -2.067951531e-37   ub1 = -1.771295037e-18 lub1 = 3.069870772e-24 wub1 = -1.925929944e-40 pub1 = -3.851859889e-46   uc1 = -5.462573950e-12 luc1 = 1.179612064e-16   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 2.75e-6   sbref = 2.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.194 pmos  lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.134757541e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.624638780e-8   k1 = 4.594670852e-01 lk1 = 2.227608917e-8   k2 = 3.309204087e-02 lk2 = 2.206364919e-9   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 1.810707000e+00 ldsub = -8.494385269e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-1.538385848e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.527858677e-8   nfactor = {3.469660796e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.448540484e-7   eta0 = -7.579850000e-02 leta0 = 3.099302733e-7   etab = -1.773594460e+00 letab = 9.715272818e-7   u0 = 8.096513985e-03 lu0 = -2.207047913e-9   ua = -4.898988585e-10 lua = -5.130754485e-16   ub = 3.687512904e-19 lub = 2.885045525e-25   uc = -9.389506674e-11 luc = 4.182499626e-17 wuc = -2.584939414e-32   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 3.593705900e+03 lvsat = 3.841069188e-2   a0 = 1.444354922e+00 la0 = -3.297923386e-7   ags = 3.137501710e-01 lags = 5.128542501e-7   a1 = 0.0   a2 = 6.137565000e-01 la2 = 1.951412832e-7   b0 = -3.703465515e-08 lb0 = 2.028665822e-14   b1 = -1.089790777e-08 lb1 = 5.969601431e-15   keta = 2.863008571e-03 lketa = -1.754711681e-8   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 7.996163666e-01 lpclm = -4.166881379e-7   pdiblc1 = 8.001533923e-01 lpdiblc1 = -4.311635851e-7   pdiblc2 = 8.716435937e-04 lpdiblc2 = -4.627431164e-10   pdiblcb = -3.618407354e-01 lpdiblcb = 1.433783016e-7   drout = 6.746922664e-01 ldrout = 1.781954438e-7   pscbe1 = 800000000.0   pscbe2 = 9.037747670e-09 lpscbe2 = 6.043307442e-17   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 5.158004358e-11 lalpha0 = 2.652324163e-17   alpha1 = -3.191100000e-10 lalpha1 = 2.295779803e-16 walpha1 = -5.169878828e-32   beta0 = 4.173312430e+00 lbeta0 = 2.187155785e-6   agidl = 1.196873537e-09 lagidl = -1.080497400e-16   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.182767825e-01 lkt1 = -4.689130247e-8   kt2 = -4.244640755e-02 lkt2 = -9.365633704e-9   at = -4.318645350e+03 lat = 4.618764596e-2   ute = -1.930957550e+00 lute = 9.653754070e-7   ua1 = -2.722113345e-09 lua1 = 2.215209410e-15 pua1 = 2.067951531e-37   ub1 = 3.302164085e-18 lub1 = -2.245972860e-24   uc1 = 2.982595129e-10 luc1 = -2.002712032e-16 puc1 = -2.584939414e-38   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.75e-6   sbref = 1.74e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.195 pmos  lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.134907458e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.632850865e-8   k1 = 8.144968549e-02 lk1 = 2.293445703e-7   k2 = 2.317871316e-01 lk2 = -1.066338384e-07 pk2 = 6.938893904e-30   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = -2.189838204e-01 ldsub = 2.623753622e-7   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-9.957617728e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.444500353e-8   nfactor = {1.608868100e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.361566913e-8   eta0 = 0.49   etab = -6.25e-6   u0 = 7.145917060e-03 lu0 = -1.686334683e-9   ua = 1.243079395e-10 lua = -8.495225773e-16   ub = -7.749310185e-19 lub = 9.149851292e-25   uc = -3.874084833e-11 luc = 1.161289427e-17   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = -1.611895310e+04 lvsat = 4.920879366e-2   a0 = 4.563589192e-01 la0 = 2.114071720e-7   ags = 1.25   a1 = 0.0   a2 = 1.586399074e+00 la2 = -3.376480027e-7   b0 = 0.0   b1 = 0.0   keta = -3.030398915e-02 lketa = 6.209353634e-10   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = -8.993470467e-01 lpclm = 5.139615458e-07 wpclm = -2.775557562e-23 ppclm = -6.938893904e-30   pdiblc1 = -1.950887668e-01 lpdiblc1 = 1.140051886e-07 wpdiblc1 = -6.938893904e-24 ppdiblc1 = -5.204170428e-30   pdiblc2 = -7.914824152e-03 lpdiblc2 = 4.350264253e-09 wpdiblc2 = -2.439454888e-25 ppdiblc2 = -1.287490080e-31   pdiblcb = 4.868147087e-02 lpdiblcb = -8.149549999e-08 ppdiblcb = -1.387778781e-29   drout = 1.002257968e+00 ldrout = -1.236858569e-9   pscbe1 = 8.000374601e+08 lpscbe1 = -2.051970354e-2   pscbe2 = 8.946288049e-09 lpscbe2 = 1.105323681e-16   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 7.071369012e+00 lbeta0 = 5.996728401e-7   agidl = -1.295214076e-09 lagidl = 1.257053552e-15   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -4.595234360e-01 lkt1 = -2.429741685e-8   kt2 = -8.004402210e-02 lkt2 = 1.122939961e-08 wkt2 = -2.775557562e-23   at = 5.017366490e+04 lat = 1.633812071e-2   ute = 1.368337730e-01 lute = -1.673089850e-07 pute = -2.775557562e-29   ua1 = 2.547029727e-09 lua1 = -6.710954362e-16   ub1 = -1.813522802e-18 lub1 = 5.562725253e-25   uc1 = -7.808557540e-11 luc1 = 5.881227590e-18   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.196 pmos  lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -2.38875e-8   vth0 = {-1.04649+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.85164386   k2 = -0.12631492   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 0.66213569   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-0.14808597+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}   nfactor = {1.7889224+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}   eta0 = 0.49   etab = -6.25e-6   u0 = 0.0014828   ua = -2.728593e-9   ub = 2.2978089e-18   uc = 2.58041e-13   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 149136.0   a0 = 1.166315   ags = 1.25   a1 = 0.0   a2 = 0.45249595   b0 = 0.0   b1 = 0.0   keta = -0.028218739   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 0.82665932   pdiblc1 = 0.18776805   pdiblc2 = 0.0066944085   pdiblcb = -0.225   drout = 0.9981043   pscbe1 = 799968550.0   pscbe2 = 9.3174823e-9   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 9.0852145   agidl = 2.9262738e-9   bgidl = 1000000000.0   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -1.46875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = -0.54112   kt2 = -0.042333   at = 105041.0   ute = -0.42503   ua1 = 2.9333e-10   ub1 = 5.4574e-20   uc1 = -5.8335e-11   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.1e-6   sbref = 1.1e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















* Well Proximity Effect Parameters





















* .model sky130_fd_pr__pfet_01v8_hvt__model.197 pmos  lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 4.2e-7   level = 54.0   version = 4.5   binunit = 2.0   mobmod = 0.0   capmod = 2.0   igcmod = 0.0   igbmod = 0.0   geomod = 0.0   diomod = 1.0   rdsmod = 0.0   rbodymod = 1.0   rgatemod = 0.0   permod = 1.0   acnqsmod = 0.0   trnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   tempmod = 0.0   toxe = {4.384395e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.0365*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}   toxm = 4.23e-9   dtox = 0.0   epsrox = 3.9   xj = 1.5e-7   ngate = 1.0e+23   ndep = 1.7e+17   nsd = 1.0e+20   rsh = 1.0   rshg = 0.1   wint = 3.1884e-8   lint = -3.23875e-8   vth0 = {-1.590239467e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.330962758e-07 wvth0 = 3.079070308e-07 pvth0 = -7.536794346e-14   k1 = -1.996351050e+00 lk1 = 6.971179541e-07 wk1 = 7.075692627e-07 pk1 = -1.731952663e-13   k2 = -2.704070119e-01 lk2 = 3.527014180e-08 wk2 = 2.357592592e-07 pk2 = -5.770797268e-14   k3 = -13.778   k3b = 2.0   w0 = 0.0   dvt0 = 4.05   dvt1 = 0.3   dvt2 = 0.03   dvt0w = -4.254   dvt1w = 1147200.0   dvt2w = -0.00896   dsub = 7.046964934e+00 ldsub = -1.562846578e-06 wdsub = -1.827541316e-06 pdsub = 4.473364257e-13   minv = 0.0   voffl = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   phin = 0.0   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   cit = 1.0e-5   voff = {-2.108998367e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.799823320e-07 wvoff = 8.014086043e-07 pvoff = -1.961647911e-13   nfactor = {4.301268408e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.009054626e-05 wnfactor = -1.492524072e-05 pnfactor = 3.653325797e-12   eta0 = 8.230920372e+00 leta0 = -1.894783784e-06 weta0 = -2.757563546e-06 peta0 = 6.749826169e-13   etab = 4.497324014e-01 letab = -1.100847784e-07 wetab = -1.586332861e-07 petab = 3.882946261e-14   u0 = 2.685845234e-02 lu0 = -6.211325302e-09 wu0 = -1.256791649e-08 pu0 = 3.076311759e-15   ua = -1.029761455e-08 lua = 1.852707249e-15 wua = 7.021962449e-16 pua = -1.718800859e-22   ub = 2.045204657e-17 lub = -4.443703525e-24 wub = -4.348982753e-24 pub = 1.064522253e-30   uc = -3.478207221e-10 luc = 8.520097923e-17 wuc = 1.735219870e-16 puc = -4.247384438e-23   ud = 0.0   up = 0.0   lp = 1.0   eu = 1.67   vtl = 0.0   xn = 3.0   vsat = 9.884931225e+05 lvsat = -2.054536397e-01 wvsat = -1.779330477e-01 pvsat = 4.355356176e-8   a0 = 2.112539359e+00 la0 = -2.316120674e-07 wa0 = 7.438728946e-08 pa0 = -1.820814878e-14   ags = 1.249999985e+00 lags = 3.619858191e-15 wags = 5.268141479e-15 pags = -1.289509388e-21   a1 = 0.0   a2 = -9.040480416e+00 la2 = 2.323643290e-06 wa2 = 2.918491330e-06 pa2 = -7.143737154e-13   b0 = 0.0   b1 = 0.0   keta = -1.586701126e+00 lketa = 3.814775263e-07 wketa = 5.271743253e-07 pketa = -1.290390955e-13   dwg = -5.722e-9   dwb = -1.7864e-8   pclm = 2.341101211e+00 lpclm = -3.706975139e-07 wpclm = -2.410278567e-08 ppclm = 5.899759362e-15   pdiblc1 = 1.411659737e-01 lpdiblc1 = 1.140702322e-08 wpdiblc1 = 7.914155401e-08 ppdiblc1 = -1.937187388e-14   pdiblc2 = 6.842249906e-02 lpdiblc2 = -1.510949337e-08 wpdiblc2 = -1.436765013e-08 ppdiblc2 = 3.516841560e-15   pdiblcb = -9.163561431e+00 lpdiblcb = 2.187936374e-06 wpdiblcb = 3.901480314e-06 ppdiblcb = -9.549848438e-13   drout = 9.845326527e-01 ldrout = 3.321999964e-09 wdrout = 5.355953903e-15 pdrout = -1.311003750e-21   pscbe1 = 1.288436647e+09 lpscbe1 = -1.195647786e+02 wpscbe1 = -1.740870784e+02 ppscbe1 = 4.261216461e-5   pscbe2 = 1.551291865e-08 lpscbe2 = -1.516487932e-15 wpscbe2 = -2.600309662e-15 ppscbe2 = 6.364907976e-22   pvag = 0.0   delta = 0.01   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   lambda = 0.0   lc = 5.0e-9   rdsw = 531.92   rsw = 0.0   rdw = 0.0   rdswmin = 0.0   rdwmin = 0.0   rswmin = 0.0   prwb = -0.32348   prwg = 0.02   wr = 1.0   alpha0 = 1.0e-10   alpha1 = 1.0e-10   beta0 = 2.401315341e+01 lbeta0 = -3.653986246e-06 wbeta0 = -3.524254723e-06 pbeta0 = 8.626494497e-13   agidl = -1.520812651e-07 lagidl = 3.794197034e-14 wagidl = 5.212415942e-14 pagidl = -1.275869112e-20   bgidl = 1.000000010e+09 lbgidl = -2.519254684e-06 wbgidl = -3.666381836e-06 pbgidl = 8.974385262e-13   cgidl = 300.0   egidl = 0.1   toxref = 4.23e-9   dlcig = 0.0   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   nigc = 1.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   vfbsdoff = 0.0   dlc = -2.31875e-8   dwc = 2.252e-8   xpart = 0.0   cgso = 6.9684e-11   cgdo = 6.9684e-11   cgbo = 0.0   cgdl = 8.82664e-12   cgsl = 8.82664e-12   clc = 1.0e-7   cle = 0.6   cf = 1.2e-11   ckappas = 0.6   vfbcv = -0.1446893   acde = 0.552   moin = 14.504   noff = 4.0   voffcv = -0.1375   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   ef = 0.88   noia = 1.2e+41   noib = 2.0e+25   noic = 0.0   em = 41000000.0   ntnoi = 1.0   lintnoi = -6.0e-8   af = 1.0   kf = 0.0   tnoia = 1.5   tnoib = 3.5   rnoia = 0.577   rnoib = 0.37   xl = 0.0   xw = 0.0   dmcg = 0.0   dmdg = 0.0   dmcgt = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   jss = 2.17e-5   jsws = 8.2e-10   ijthsfwd = 0.1   ijthsrev = 0.1   bvs = 12.8   xjbvs = 1.0   pbs = 0.6587   cjs = 0.000792710451   mjs = 0.34629   pbsws = 0.7418   cjsws = 1.01401195e-10   mjsws = 0.26859   pbswgs = 1.3925   cjswgs = 2.7096997e-10   mjswgs = 0.70393   tnom = 30.0   kt1 = 5.950906407e-01 lkt1 = -2.781159596e-07 wkt1 = -4.531597434e-07 pkt1 = 1.109221762e-13   kt2 = 1.131083619e+00 lkt2 = -2.872230530e-07 wkt2 = -4.015742596e-07 pkt2 = 9.829533938e-14   at = 1.185891568e+05 lat = -3.316250091e-03 wat = 1.683177773e-01 pat = -4.119998395e-8   ute = -2.299514599e+00 lute = 4.588269676e-07 wute = -3.451785524e-15 pute = 8.449108080e-22   ua1 = -1.102559745e-09 lua1 = 3.416789124e-16 wua1 = -9.065908965e-16 pua1 = 2.219107867e-22   ub1 = 5.406746700e-18 lub1 = -1.310078073e-24 wub1 = -1.620301706e-25 pub1 = 3.966093500e-32   uc1 = -9.345371040e-10 luc1 = 2.144723700e-16 wuc1 = 3.744968574e-16 puc1 = -9.166746826e-23   kt1l = 0.0   prt = 0.0   tvoff = 0.0   njs = 1.2556   tpb = 0.0019551   tcj = 0.0012407   tpbsw = 0.00014242   tcjsw = 0.0   tpbswg = 0.0   tcjswg = 2.0e-12   xtis = 2.0   tvfbsdoff = 0.0   ll = 0.0   wl = 0.0   lln = 1.0   wln = 1.0   lw = 0.0   ww = 0.0   lwn = 1.0   wwn = 1.0   lwl = 0.0   wwl = 0.0   llc = 0.0   wlc = 0.0   lwc = 0.0   wwc = 0.0   lwlc = 0.0   wwlc = 0.0   saref = 1.04e-6   sbref = 1.04e-6   kvth0 = 2.65e-8   lkvth0 = 0.0   wkvth0 = 2.5e-7   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   wlod = 0.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = 4.5e-8   lku0 = 0.0   wku0 = 2.5e-7   pku0 = 0.0   tku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = 0.4   steta0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* Model Flag Parameters
* Process Parameters



















* Basic Model Parameters










* Parameters FOR Asymmetric AND Bias-Dependent RDS Model


































































* Impact Ionization Current Model Parameters









* Gidl Induced Drain Leakage Model Parameters



* Gate Dielectric Tunneling Current Model Parameters




* Charge AND Capacitance Model Parameters






















* High-Speed/RF Model Parameters

















* Flicker AND Thermal Noise Model Parameters








* Layout-Dependent Parasitics Model Parameters













* Asymmetric Source/Drain Junction Diode Model Parameters








* Temperature Dependence Parameters















* DW AND DL Parameters




















* Stress Parameters
















.ENDS sky130_fd_pr__pfet_01v8_hvt





















* Well Proximity Effect Parameters
