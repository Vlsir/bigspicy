** Translated using xdm 2.6.0 on Nov_14_2022_16_05_19_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 52
.PARAM 
+ SKY130_FD_PR__PFET_01V8__AJUNCTION_MULT=0.93001 SKY130_FD_PR__PFET_01V8__PJUNCTION_MULT=0.93439
.INCLUDE sky130_fd_pr__pfet_01v8__ff.pm3.spice

