** Translated using xdm 2.6.0 on Nov_14_2022_16_05_17_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_G5V0D10V5__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_G5V0D10V5__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_G5V0D10V5__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_G5V0D10V5__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__nfet_g5v0d10v5 d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__nfet_g5v0d10v5 d g s b sky130_fd_pr__nfet_g5v0d10v5__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__nfet_g5v0d10v5__model.0 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.1 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.2 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.778154642625+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.87586169956661e-8   k1 = 0.88325   k2 = -0.042248784952 lk2 = 1.16867712579414e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110512.045 lvsat = -0.03824205254562   ua = -1.020396686767e-10 lua = 3.35813406336751e-16   ub = 1.57307850057e-18 lub = 9.27522742441469e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.040631002942 lu0 = 1.04171351134268e-8   a0 = 1.0357342704916 la0 = -7.52545466177932e-7   keta = -0.017231666883 lketa = -3.22227534749394e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1458383692056 lags = 8.00146113822516e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05983857844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.37183144701528e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.25924117019 lpclm = 5.89615966148369e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4769366 lbeta0 = 1.98858673237224e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414374908 lkt1 = 9.17809261094877e-8   kt2 = -0.019151   at = 237632.72 lat = -0.61187284072992   ute = -1.33741636 lute = 3.05936420364959e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.3 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793057696002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.08961150241902e-9   k1 = 0.88325   k2 = -0.0433694140834 lk2 = 1.60366456370324e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93650.9059 lvsat = 0.0272067519859476   ua = 1.078566180374e-10 lua = -4.78927576439021e-16 wua = -9.86076131526265e-32 pua = -5.64237288394698e-37   ub = 1.557827562126e-18 lub = 9.86721334139483e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04291014826 lu0 = 1.57032259784664e-9   a0 = 0.464123513818 la0 = 1.46623942491356e-6   keta = -0.039525786114 lketa = 5.43149023204025e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.124583717364 lags = 1.62517433138072e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.99638655686+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.90885493463824e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60454395626 lpclm = -7.50723759161242e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.807652176 lbeta0 = 1.08388778381601e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284642e-8   kt2 = -0.019151   at = 140212.352 lat = -0.233722433167872   ute = -1.22096728 lute = -1.4607652072992e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.4 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.767943200548+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.81667272656634e-8   k1 = 0.88325   k2 = -0.0416548695192 lk2 = 1.28104968614294e-08 wk2 = -2.11758236813575e-22   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 120367.385308 lvsat = -0.0230639374614039   ua = -1.423282782092e-10 lua = -8.17066900515378e-18   ub = 1.764175457908e-18 lub = 5.98449704911823e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0423086912832 lu0 = 2.70204569784469e-9   a0 = 1.751557912936 la0 = -9.56243488105244e-7   keta = 0.00389404708800001 lketa = -2.7385418946476e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.111605965704 lags = 1.86936837860588e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.89703829368+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.9482249268604e-9   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.09229740672 lpclm = 2.13137789329006e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 26.983043248 lbeta0 = 4.86394768300626e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.38154636 lkt1 = 1.65891803649599e-8   kt2 = -0.019151   at = 8946.91199999999 lat = 0.013271344291968   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.0171671272e-18 lub1 = 4.98007194556099e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.5 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.77380195906+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.30014348461777e-8   k1 = 0.88325   k2 = -0.037465940574 lk2 = 9.11738630189907e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 52828.968256 lvsat = 0.0364803623946532   ua = -1.65085135622e-10 lua = 1.18925957368376e-17   ub = 2.9580482434e-18 lub = -4.54111522198202e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04676425556352 lu0 = -1.22614017199951e-9   a0 = -0.88469447588 la0 = 1.36797152296094e-6   keta = -0.08343023544 lketa = 4.96028122043799e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.8805025302 lags = -4.90950053675407e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.978786954+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.60207868167443e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.030374875 lpclm = 2.0845620890955e-06 ppclm = -3.23117426778526e-27   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.60713526000001e-06 lalpha0 = 8.69281170991464e-12   alpha1 = 0.0   beta0 = 22.33680724 lbeta0 = 8.96023661215535e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.33546456 lkt1 = -2.40381934598401e-8   kt2 = -0.019151   at = 6959.10000000001 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397719e-7   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -1.0286723354e-17 lub1 = 6.02547366812715e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.6 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.75996795518+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.24311899149256e-8   k1 = 0.88325   k2 = -0.019352346668 lk2 = -3.22949139381116e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93236.223172 lvsat = 0.0089373227827306   ua = -3.14415783446e-10 lua = 1.13681741196998e-16   ub = 1.4486398548e-18 lub = 5.74755574173547e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03972026583648 lu0 = 3.57529680958113e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.9960013028+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.77547066753809e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.032134724 lpclm = -2.95470392846365e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.66616278e-05 lalpha0 = 4.76035632919197e-13   alpha1 = 0.0   beta0 = 31.92270996 lbeta0 = 2.42614022570544e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10799999999 lat = 0.015430120515312   ute = -1.12187464 lute = -8.535811348896e-8   ua1 = 2.0117e-9   ub1 = -1.687818e-18 lub1 = 1.64150218248e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.7 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.684534974+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.87624292385363e-8   k1 = 0.88325   k2 = -0.00719142434 lk2 = -9.08662938017976e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 43946.678464 lvsat = 0.0326769419377129   ua = 2.78994770932e-10 lua = -1.72126144571405e-16   ub = -2.01261184512e-17 lub = 1.09659358656422e-23   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.00318094097999999 lu0 = 2.11739510761567e-8   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.309048226400001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.43106625229609e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.0383260320000005 lpclm = 4.75699339251648e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.979747388e-05 lalpha0 = -5.85066072966768e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4470572 lkt1 = 3.67619272992e-8   kt2 = -0.019151   at = -4343.23199999999 lat = 0.020586679287552   ute = -1.30100818 lute = 9.19048182479615e-10   ua1 = -1.776800572e-09 lua1 = 1.82467826149579e-15   ub1 = 6.49752798e-18 lub1 = -3.77820707817528e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.8 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.9 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.10 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.778154642625+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.87586169956653e-8   k1 = 0.88325   k2 = -0.042248784952 lk2 = 1.16867712579414e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110512.045 lvsat = -0.0382420525456202   ua = -1.020396686767e-10 lua = 3.35813406336751e-16   ub = 1.57307850057e-18 lub = 9.27522742441478e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0406310029420001 lu0 = 1.04171351134272e-8   a0 = 1.0357342704916 la0 = -7.52545466177935e-7   keta = -0.017231666883 lketa = -3.22227534749394e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1458383692056 lags = 8.00146113822522e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05983857844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.37183144701522e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.25924117019 lpclm = 5.89615966148368e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4769366 lbeta0 = 1.98858673237224e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414374908 lkt1 = 9.17809261094885e-8   kt2 = -0.019151   at = 237632.72 lat = -0.61187284072992   ute = -1.33741636 lute = 3.05936420364954e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.11 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793057696001999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.0896115024186e-9   k1 = 0.88325   k2 = -0.0433694140834 lk2 = 1.60366456370325e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93650.9059 lvsat = 0.0272067519859474   ua = 1.078566180374e-10 lua = -4.78927576439022e-16 pua = -2.25694915357879e-36   ub = 1.557827562126e-18 lub = 9.86721334139476e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04291014826 lu0 = 1.57032259784658e-9   a0 = 0.464123513817999 la0 = 1.46623942491356e-6   keta = -0.039525786114 lketa = 5.43149023204026e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.124583717364 lags = 1.62517433138073e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.99638655686+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.90885493463823e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60454395626 lpclm = -7.50723759161242e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.807652176 lbeta0 = 1.08388778381601e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284635e-8   kt2 = -0.019151   at = 140212.352 lat = -0.233722433167872   ute = -1.22096728 lute = -1.46076520729919e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.12 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.770789820952902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.28104238334653e-08 wvth0 = -5.66277001566508e-08 pvth0 = 1.06552719211959e-13   k1 = 0.88325   k2 = -0.0417969379360867 lk2 = 1.30778179091064e-08 wk2 = 2.82616105025333e-09 pk2 = -5.31780637395508e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 128245.486059573 lvsat = -0.0378876554471903 wvsat = -0.156718727370807 pvsat = 2.94887599295094e-7   ua = -1.42366880902883e-10 lua = -8.09803278702333e-18 wua = 7.67921764117603e-19 pua = -1.44494923654526e-24   ub = 1.38681443190766e-18 lub = 1.30850579643099e-24 wub = 7.50682704106159e-24 pub = -1.41251160062349e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419476116654196 lu0 = 3.38146610552653e-09 wu0 = 7.18294167116219e-09 pu0 = -1.35156816343581e-14   a0 = 1.73734581918016 la0 = -9.29501500858886e-07 wa0 = 2.82720584176931e-07 pa0 = -5.31977229128352e-13   keta = 0.00389404708799999 lketa = -2.7385418946476e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.134951404264494 lags = 1.43009220229375e-07 wags = -4.64409828775491e-07 pags = 8.73850252577796e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.889081411920912+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.10237302387844e-08 wnfactor = 1.5828591464452e-07 pnfactor = -2.97836475288047e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.09229740672 lpclm = 2.13137789329006e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 27.0486940875965 lbeta0 = 4.74041669979141e-06 wbeta0 = -1.30598939475672e-06 pbeta0 = 2.45739666079223e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.38154636 lkt1 = 1.65891803649599e-8   kt2 = -0.019151   at = 8946.91200000001 lat = 0.013271344291968   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.0171671272e-18 lub1 = 4.980071945561e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.13 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.759568857035493+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.27032295777554e-08 wvth0 = 2.83138500783254e-07 pvth0 = -1.92997395119899e-13   k1 = 0.88325   k2 = -0.0367555984895665 lk2 = 8.63319156483415e-09 wk2 = -1.41308052512675e-08 pk2 = 9.63206556825342e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 13438.4644981362 lvsat = 0.0633303478141485 wvsat = 0.783593636854029 pvsat = -5.34125632250634e-7   ua = -1.64892122153586e-10 lua = 1.17610308082825e-17 wua = -3.83960882057855e-18 pua = 2.61721559802516e-24   ub = 4.84485337340168e-18 lub = -1.74022582379202e-24 wub = -3.7534135205308e-23 pub = 2.55846177848054e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0485696536524221 lu0 = -2.45676450372631e-09 wu0 = -3.59147083558093e-08 pu0 = 2.44807581448197e-14   a0 = -0.813634007100815 la0 = 1.31953414926417e-06 wa0 = -1.41360292088465e-06 pa0 = 9.63562640580134e-13   keta = -0.08343023544 lketa = 4.96028122043798e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.763775337397529 lags = -4.11384596882302e-07 wags = 2.32204914387745e-06 pags = -1.58279229023604e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.01857136279544+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.03139272090433e-07 wnfactor = -7.91429573222574e-07 pnfactor = 5.39466888573125e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.030374875 lpclm = 2.0845620890955e-06 ppclm = 1.29246970711411e-26   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.60713525999998e-06 lalpha0 = 8.69281170991463e-12   alpha1 = 0.0   beta0 = 22.0085530420179 lbeta0 = 9.18398649065111e-06 wbeta0 = 6.52994697378402e-06 pbeta0 = -4.45104693542181e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.33546456 lkt1 = -2.40381934598398e-8   kt2 = -0.019151   at = 6959.10000000003 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397724e-7   ua1 = 6.387700286e-09 lua1 = -2.98283933094789e-15   ub1 = -1.0286723354e-17 lub1 = 6.02547366812714e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.14 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.75996795518+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.24311899149262e-8   k1 = 0.88325   k2 = -0.019352346668 lk2 = -3.22949139381115e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93236.2231720001 lvsat = 0.00893732278273063   ua = -3.14415783446e-10 lua = 1.13681741196998e-16   ub = 1.4486398548e-18 lub = 5.74755574173548e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03972026583648 lu0 = 3.57529680958114e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.9960013028+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.77547066753809e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.032134724 lpclm = -2.95470392846365e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.66616278e-05 lalpha0 = 4.76035632919197e-13   alpha1 = 0.0   beta0 = 31.92270996 lbeta0 = 2.42614022570543e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000007 lat = 0.0154301205153121   ute = -1.12187464 lute = -8.535811348896e-8   ua1 = 2.0117e-9   ub1 = -1.687818e-18 lub1 = 1.64150218248e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.15 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.625583752529145+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.07155459742872e-07 wvth0 = 1.17271417276842e-06 pvth0 = -5.6482136331549e-13   k1 = 0.88325   k2 = -0.0252814694323099 lk2 = -3.73812422100003e-10 wk2 = 3.59864507239426e-07 pk2 = -1.73323701808769e-13   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -125620.496754038 lvsat = 0.114346597941028 wvsat = 3.37319269479107 pvsat = -1.62465103674839e-6   ua = 6.30267207424107e-10 lua = -3.41311595793717e-16 wua = -6.98784782569516e-15 pua = 3.36559907537652e-21   ub = -6.30425167429598e-17 lub = 3.16360182732922e-23 wub = 8.53734108729249e-22 pub = -4.11189081191921e-28   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = -0.0518803637944942 lu0 = 4.7693457662525e-08 wu0 = 1.09533222330422e-06 pu0 = -5.27551430703349e-13   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {-0.34878192911839+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.59941310012866e-07 wnfactor = 1.30861876548608e-05 pnfactor = -6.30277907733656e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.29880685161122 lpclm = 1.60134667278262e-06 wpclm = 4.6492486294097e-05 ppclm = -2.23924551287437e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.979747388e-05 lalpha0 = -5.85066072966765e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4470572 lkt1 = 3.67619272992003e-8   kt2 = -0.019151   at = -94554.742526939 lat = 0.0640357903717049 wat = 1.79457379002896 pat = -8.64331341934387e-7   ute = -1.30100818 lute = 9.19048182478768e-10   ua1 = -1.77680057199999e-09 lua1 = 1.82467826149579e-15   ub1 = 2.5189457364984e-18 lub1 = -1.86197864074414e-24 wub1 = 7.91457694695229e-23 pub1 = -3.81194518242232e-29   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.16 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.17 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.18 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.778154642625+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.87586169956653e-8   k1 = 0.88325   k2 = -0.042248784952 lk2 = 1.16867712579414e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110512.045 lvsat = -0.0382420525456197   ua = -1.020396686767e-10 lua = 3.35813406336751e-16   ub = 1.57307850057e-18 lub = 9.2752274244146e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.040631002942 lu0 = 1.0417135113427e-8   a0 = 1.0357342704916 la0 = -7.52545466177932e-7   keta = -0.017231666883 lketa = -3.22227534749394e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1458383692056 lags = 8.00146113822518e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05983857844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.37183144701528e-07 wnfactor = -6.7762635780344e-21   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.25924117019 lpclm = 5.89615966148369e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4769366 lbeta0 = 1.98858673237225e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414374908 lkt1 = 9.17809261094885e-8   kt2 = -0.019151   at = 237632.72 lat = -0.61187284072992   ute = -1.33741636 lute = 3.05936420364964e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.19 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793057696002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.0896115024186e-9   k1 = 0.88325   k2 = -0.0433694140834 lk2 = 1.60366456370324e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93650.9058999999 lvsat = 0.0272067519859478   ua = 1.078566180374e-10 lua = -4.78927576439021e-16 wua = 9.86076131526265e-32 pua = 9.4039548065783e-37   ub = 1.557827562126e-18 lub = 9.86721334139482e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04291014826 lu0 = 1.57032259784664e-9   a0 = 0.464123513818 la0 = 1.46623942491356e-6   keta = -0.039525786114 lketa = 5.43149023204026e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.124583717364 lags = 1.62517433138072e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.99638655686+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.90885493463822e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60454395626 lpclm = -7.50723759161242e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.807652176 lbeta0 = 1.083887783816e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284644e-8   kt2 = -0.019151   at = 140212.352 lat = -0.233722433167872   ute = -1.22096728 lute = -1.46076520729919e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.20 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.756214107646096+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.02366107172314e-08 wvth0 = 1.60447785941653e-07 pvth0 = -3.01904330148109e-13   k1 = 0.88325   k2 = -0.0387547340824761 lk2 = 7.35349761881392e-09 wk2 = -4.24812531690077e-08 pk2 = 7.99342552879194e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 125089.068304631 lvsat = -0.0319484261684519 wvsat = -0.109710330315998 pvsat = 2.06434907094474e-7   ua = -1.39591842544251e-10 lua = -1.33196448640064e-17 wua = -4.05606079593785e-17 pua = 7.6320300118254e-23   ub = 1.45747620459133e-18 lub = 1.17554606112559e-24 wub = 6.45446422827822e-24 pub = -1.21449522526405e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0424421793482145 lu0 = 2.45086974914304e-09 wu0 = -1.82634056860387e-10 pu0 = 3.43650816214475e-16   a0 = 2.74604469532612 la0 = -2.82750561937466e-06 wa0 = -1.4739789412912e-05 pa0 = 2.77349183917541e-11   keta = 0.0326905624023213 lketa = -8.15699788364542e-08 wketa = -4.28865293122543e-07 pketa = 8.0696837468993e-13   a1 = 0.0   a2 = 0.65972622   ags = -0.0439211997733036 lags = 4.7958235140064e-07 wags = 2.19953235051006e-06 pags = -4.13871925388435e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.859623394282952+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.64529967150028e-08 wnfactor = 5.97002934089903e-07 pnfactor = -1.12334221288918e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.764658011442073 lpclm = -1.05200012949782e-06 wpclm = -1.00134382469804e-05 ppclm = 1.88416458892953e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.24487319954767e-05 lalpha0 = 3.79764573495911e-12 walpha0 = 3.00579806241085e-11 palpha0 = -5.6558178429625e-17   alpha1 = 0.0   beta0 = 27.4407116835608 lbeta0 = 4.00278227859132e-06 wbeta0 = -7.14429098671557e-06 pbeta0 = 1.34429551150794e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.398990335838576 lkt1 = 4.94123932859548e-08 wkt1 = 2.59792399516929e-07 pkt1 = -4.88834731457432e-13   kt2 = -0.019151   at = 8946.912 lat = 0.013271344291968   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.54083528187405e-18 lub1 = 1.48336004644436e-24 wub1 = 7.79896783349816e-24 pub1 = -1.46748186383521e-29   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.21 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.832447423569521+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.97342500023521e-09 wvth0 = -8.02238929708263e-07 pvth0 = 5.46834935090623e-13   k1 = 0.88325   k2 = -0.0519666177576197 lk2 = 1.90015698946329e-08 wk2 = 2.12406265845039e-07 pk2 = -1.44783757425549e-13   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 29220.5532728469 lvsat = 0.0525727079501097 wvsat = 0.54855165157999 pvsat = -3.73912553576378e-7   ua = -1.78767313946746e-10 lua = 2.12188610414047e-17 wua = 2.02803039796895e-16 pua = -1.38237852834996e-22   ub = 4.49154450998334e-18 lub = -1.49939778336701e-24 wub = -3.2272321141391e-23 pub = 2.19979758935332e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0460968152384473 lu0 = -7.71188818578352e-10 wu0 = 9.13170284301934e-10 pu0 = -6.22449739910517e-16   a0 = -5.85712838783059 la0 = 4.75736148496729e-06 wa0 = 7.36989470645599e-05 pa0 = -5.02358554812983e-11   keta = -0.227412812011606 lketa = 1.47746519768343e-07 wketa = 2.14432646561271e-06 pketa = -1.46165011471439e-12   a1 = 0.0   a2 = 0.65972622   ags = 1.65813835758652 lags = -1.02101462851184e-06 wags = -1.09976617525503e-05 pags = 7.49640216636138e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.16586145098524+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.03537498643775e-07 wnfactor = -2.98501467044949e-06 pnfactor = 2.03469345990651e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -5.39217789861036 lpclm = 4.37608805489717e-06 wpclm = 5.00671912349021e-05 ppclm = -3.41275999645937e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.46984752826162e-05 lalpha0 = 1.81419106225862e-12 walpha0 = -1.50289903120542e-10 palpha0 = 1.02443008403474e-16   alpha1 = 0.0   beta0 = 20.0484650621958 lbeta0 = 1.05200530208651e-05 wbeta0 = 3.57214549335776e-05 pbeta0 = -2.4349029655104e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.24824468080712 lkt1 = -8.3490403033358e-08 wkt1 = -1.29896199758463e-06 pkt1 = 8.85419260185598e-13   kt2 = -0.019151   at = 6959.09999999992 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397719e-7   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -7.66838258062975e-18 lub1 = 4.24071833673014e-24 wub1 = -3.89948391674907e-23 pub1 = 2.65802861907717e-29   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.22 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.75996795518+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.24311899149254e-8   k1 = 0.88325   k2 = -0.019352346668 lk2 = -3.22949139381116e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93236.2231719998 lvsat = 0.00893732278273074   ua = -3.14415783446e-10 lua = 1.13681741196998e-16   ub = 1.4486398548e-18 lub = 5.74755574173547e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0397202658364799 lu0 = 3.57529680958114e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.996001302799998+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.77547066753801e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.032134724 lpclm = -2.95470392846365e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.66616278e-05 lalpha0 = 4.76035632919197e-13   alpha1 = 0.0   beta0 = 31.92270996 lbeta0 = 2.42614022570546e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000001 lat = 0.015430120515312   ute = -1.12187464 lute = -8.53581134889591e-8   ua1 = 2.0117e-9   ub1 = -1.687818e-18 lub1 = 1.64150218248e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.23 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.760747822249842+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.20555778588771e-08 wvth0 = -8.40278640690964e-07 pvth0 = 4.04708443387837e-13   k1 = 0.88325   k2 = -0.00554221038762165 lk2 = -9.88095019134748e-09 wk2 = 6.5888551335764e-08 pk2 = -3.1734298311152e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 96967.6688525372 lvsat = 0.00714012421093946 wvsat = 0.0581964931153074 pvsat = -2.80295261580845e-8   ua = 4.77397221697866e-11 lua = -6.07453879057675e-17 wua = 1.68770954604305e-15 pua = -8.12861674917992e-22   ub = -9.19507662186424e-18 lub = 5.70115260312821e-24 wub = 5.17864445982586e-23 pub = -2.49422160305268e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0162714233023377 lu0 = 1.48691035323554e-08 wu0 = 8.03505204461579e-08 pu0 = -3.86997032656057e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.848251891674366+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.65932712984739e-08 wnfactor = -4.74118676278518e-06 pnfactor = 2.28352622768081e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.37545891561123 lpclm = -6.49947994279328e-07 wpclm = -2.31211574579847e-05 ppclm = 1.11359817934339e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.979747388e-05 lalpha0 = -5.85066072966767e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.447057200000001 lkt1 = 3.67619272991999e-8   kt2 = -0.019151   at = 85868.2785269392 lat = -0.0228624317966008 wat = -0.892458684759566 pat = 4.29840231092858e-7   ute = -1.30100818 lute = 9.19048182479615e-10   ua1 = -1.77680057199999e-09 lua1 = 1.82467826149579e-15   ub1 = 7.83325397999999e-18 lub1 = -4.42154080591128e-24 wub1 = 2.35098870164458e-38   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.24 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.25 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.784341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.040766   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 105660.0   ua = -5.94326e-11   ub = 1.69076e-18   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0419527   a0 = 0.9402534   keta = -0.02132   a1 = 0.0   a2 = 0.65972622   ags = 0.1559904   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00437+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.33405   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 24.0   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 160000.0   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.26 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.778154642625001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.87586169956653e-8   k1 = 0.88325   k2 = -0.042248784952 lk2 = 1.16867712579412e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 110512.045 lvsat = -0.0382420525456197   ua = -1.020396686767e-10 lua = 3.35813406336751e-16   ub = 1.57307850057e-18 lub = 9.2752274244146e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.040631002942 lu0 = 1.0417135113427e-8   a0 = 1.0357342704916 la0 = -7.52545466177935e-7   keta = -0.017231666883 lketa = -3.22227534749395e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1458383692056 lags = 8.00146113822514e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05983857844+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.37183144701525e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.25924117019 lpclm = 5.89615966148368e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.4769366 lbeta0 = 1.98858673237225e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414374908 lkt1 = 9.17809261094885e-8   kt2 = -0.019151   at = 237632.72 lat = -0.61187284072992 wat = 8.88178419700125e-16   ute = -1.33741636 lute = 3.05936420364961e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.27 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793057696002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.0896115024186e-9   k1 = 0.88325   k2 = -0.0433694140833999 lk2 = 1.60366456370324e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93650.9059 lvsat = 0.0272067519859476   ua = 1.078566180374e-10 lua = -4.78927576439022e-16 wua = -9.86076131526265e-32 pua = 5.64237288394698e-37   ub = 1.557827562126e-18 lub = 9.86721334139482e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04291014826 lu0 = 1.57032259784658e-9   a0 = 0.464123513817999 la0 = 1.46623942491355e-6   keta = -0.039525786114 lketa = 5.43149023204025e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.124583717364 lags = 1.62517433138073e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.996386556859999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.90885493463825e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.60454395626 lpclm = -7.50723759161242e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 23.807652176 lbeta0 = 1.083887783816e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284644e-8   kt2 = -0.019151   at = 140212.352 lat = -0.233722433167872   ute = -1.22096728 lute = -1.46076520729921e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.28 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.77243249106+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.97195166238262e-8   k1 = 0.88325   k2 = -0.0430488241988 lk2 = 1.54334121689332e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 113999.32848 lvsat = -0.0110815724837933   ua = -1.4369178999772e-10 lua = -5.60503613745017e-18   ub = 2.1099063704e-18 lub = -5.20900263459752e-26   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04242371833212 lu0 = 2.48560666162301e-9   a0 = 1.25611727292 la0 = -2.4004543988098e-8   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.178411933604 lags = 6.12323236451039e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.919969646040001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.70966830561209e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.24752037312 lpclm = 8.52551157316024e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.5487052852e-05 lalpha0 = -1.91936816822587e-12   alpha1 = 0.0   beta0 = 26.718552448 lbeta0 = 5.36162309395507e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 8946.912 lat = 0.013271344291968   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.29 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.751355506500001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.8301744983365e-8   k1 = 0.88325   k2 = -0.030496167176 lk2 = 4.36653784197994e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 84669.2523960001 lvsat = 0.0147768784746001   ua = -1.582675766794e-10 lua = 7.24550212943938e-18   ub = 1.22939368094001e-18 lub = 7.24201659138784e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0461891203189201 lu0 = -8.34107284411386e-10   a0 = 1.5925087242 la0 = -3.20579357528789e-7   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.5464726907 lags = -2.63263289997985e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.864130192199999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.13338966956032e-9   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.3312859758 lpclm = 9.26401928200408e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -4.93128999999983e-07 lalpha0 = 1.2169335439044e-11   alpha1 = 0.0   beta0 = 23.65926124 lbeta0 = 8.05880435741138e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.379546360000001 lkt1 = 6.00954836496017e-9   kt2 = -0.019151   at = 6959.10000000003 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397719e-7   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -1.161005899e-17 lub1 = 6.92750687770765e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.30 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.75996795518+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.24311899149254e-8   k1 = 0.88325   k2 = -0.019352346668 lk2 = -3.22949139381118e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93236.2231720001 lvsat = 0.00893732278273063   ua = -3.14415783446e-10 lua = 1.13681741196998e-16   ub = 1.4486398548e-18 lub = 5.74755574173545e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03972026583648 lu0 = 3.57529680958109e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.996001302800002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.77547066753809e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.032134724 lpclm = -2.95470392846449e-9   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.66616278e-05 lalpha0 = 4.76035632919197e-13   alpha1 = 0.0   beta0 = 31.92270996 lbeta0 = 2.42614022570546e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000001 lat = 0.015430120515312   ute = -1.12187464 lute = -8.535811348896e-8   ua1 = 2.0117e-9   ub1 = -1.687818e-18 lub1 = 1.64150218248e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.31 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.484478401510453+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.75116876586111e-07 wvth0 = 1.89284313536812e-06 pvth0 = -9.11661396346165e-13   k1 = 0.88325   k2 = 0.0288789308493381 lk2 = -2.64594109721519e-08 wk2 = -2.74638353233547e-07 pk2 = 1.32275717897993e-13   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93699.3031527703 lvsat = 0.00871428679311248 wvsat = 0.0905302977117408 pvsat = -4.36026504686921e-8   ua = 2.78903562012292e-10 lua = -1.72082215072152e-16 wua = -5.9918461263758e-16 pua = 2.88588880092314e-22   ub = -1.14234139352201e-17 lub = 6.77440007338365e-24 wub = 7.38312920491206e-23 pub = -3.55598081773702e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.00873169376153238 lu0 = 1.85005087094706e-08 wu0 = 1.54940748124702e-07 pu0 = -7.46250421637893e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.00396352110013609+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.90046402351416e-07 wnfactor = 3.61132262719409e-06 pnfactor = -1.73934298487125e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.0383260320000041 lpclm = 4.75699339251648e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.979747388e-05 lalpha0 = -5.85066072966767e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.447057200000001 lkt1 = 3.67619272991999e-8   kt2 = -0.019151   at = -88522.461417216 lat = 0.0611304266271423 wat = 0.832781581096882 pat = -4.01097589593178e-7   ute = -1.30100818 lute = 9.19048182478768e-10   ua1 = -1.776800572e-09 lua1 = 1.82467826149579e-15   ub1 = 9.58698792619199e-18 lub1 = -5.26620220881941e-24 wub1 = -1.73496162728517e-23 pub1 = 8.35619978319121e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.32 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.771046833114+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 9.16361339901898e-8   k1 = 0.88325   k2 = -0.040812483101 wk2 = 3.2040606290282e-10   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 119042.24013 wvsat = -0.0922432191620044   ua = -3.735064364141e-10 wua = 2.16489776330126e-15   ub = 2.10431281016e-18 wub = -2.85060215121485e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0409131910729 wu0 = 7.16529137512526e-9   a0 = 1.2253584785751 wa0 = -1.96521733220486e-6   keta = -0.017085144851 wketa = -2.91906786781408e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1693564933686 wags = -9.21319202138382e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.961703406239999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.94099038790746e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.64927881915 wpclm = -2.17285901079055e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.3668207519e-05 walpha0 = -6.34235369777512e-11   alpha1 = 0.0   beta0 = 26.654429715 wbeta0 = -1.8296872539447e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 179571.832 wat = -0.134907815959056   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.33 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.771046833113999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 9.16361339901898e-8   k1 = 0.88325   k2 = -0.040812483101 wk2 = 3.20406062902926e-10   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 119042.24013 wvsat = -0.0922432191620048   ua = -3.735064364141e-10 wua = 2.16489776330126e-15   ub = 2.10431281016e-18 wub = -2.85060215121486e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0409131910729 wu0 = 7.16529137512516e-9   a0 = 1.2253584785751 wa0 = -1.96521733220487e-6   keta = -0.017085144851 wketa = -2.91906786781409e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.1693564933686 wags = -9.21319202138387e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.96170340624+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.94099038790743e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.64927881915 wpclm = -2.17285901079055e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.3668207519e-05 walpha0 = -6.34235369777512e-11   alpha1 = 0.0   beta0 = 26.654429715 wbeta0 = -1.82968725394471e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 179571.832 wat = -0.134907815959056   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.34 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.756544055143592+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.14305616951575e-07 wvth0 = 1.48960871864672e-07 pvth0 = -4.51812717722111e-13   k1 = 0.88325   k2 = -0.0451417962556533 lk2 = 3.4122070414989e-08 wk2 = 1.99414054096075e-08 pk2 = -1.54645574806963e-13   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 142008.555510521 lvsat = -0.181012138090467 wvsat = -0.21710412409558 pvsat = 9.84108203317042e-7   ua = -5.2121781978952e-10 lua = 1.16420735682151e-15 wua = 2.88937739013832e-15 pua = -5.71008470814553e-21   ub = 2.10372119476241e-18 lub = 4.66289721580153e-27 wub = -3.65769780407514e-24 pub = 6.36123415302701e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0389317357267288 lu0 = 1.5617109788776e-08 wu0 = 1.17129775456419e-08 pu0 = -3.58432070382442e-14   a0 = 1.54009063173444 la0 = -2.48060426869815e-06 wa0 = -3.4765072150797e-06 pa0 = 1.19114367473021e-11   keta = -0.00299479061825494 lketa = -1.11055043173556e-07 wketa = -9.81341901440845e-08 pketa = 5.43387661936396e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.185930489753974 lags = -1.30630206574836e-07 wags = -2.76353303070881e-07 pags = 1.45196588309584e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.968954313457408+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.71490113573741e-08 wnfactor = 6.26461421385879e-07 pnfactor = -2.61955931970766e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.391451758195261 lpclm = 2.03209904539507e-06 wpclm = -9.11322030275567e-07 ppclm = -9.94297528095816e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.53439587288823e-05 lalpha0 = -9.2024021062852e-11 walpha0 = -1.43903999685919e-10 palpha0 = 6.34317712177354e-16   alpha1 = 0.0   beta0 = 26.7333637379425 lbeta0 = -6.22129236848038e-07 wbeta0 = -3.62323314918975e-05 pbeta0 = 1.41360758956157e-10   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414374908 lkt1 = 9.17809261094885e-8   kt2 = -0.019151   at = 276197.233919288 lat = -0.761566246281529 wat = -0.265823574736068 pat = 1.03183035734421e-6   ute = -1.33741636 lute = 3.05936420364961e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.35 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.797563327887086+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.49162688233909e-08 wvth0 = -3.10571313473589e-08 pvth0 = 2.46951644193847e-13   k1 = 0.88325   k2 = -0.0392477113844755 lk2 = 1.12433783919699e-08 wk2 = -2.84107235921735e-08 pk2 = 3.30397898029919e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 72899.1445155962 lvsat = 0.0872454395662283 wvsat = 0.143041019648718 pvsat = -4.13844151865997e-7   ua = 1.24759321613816e-10 lua = -1.34324077042677e-15 wua = -1.16509625838685e-16 pua = 5.9576745450034e-21   ub = 1.27804077429445e-18 lub = 3.20965374179937e-24 wub = 1.9285585774778e-24 pub = -1.53225797228385e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0437075991708213 lu0 = -2.92105368689802e-09 wu0 = -5.49679563535297e-09 pu0 = 3.09588680929396e-14   a0 = 0.265373267970066 la0 = 2.46738454031474e-06 wa0 = 1.36997709711949e-06 pa0 = -6.9008512323655e-12   keta = -0.0513107452449182 lketa = 7.6489905679667e-08 wketa = 8.12332283211357e-08 pketa = -1.52851366805269e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.10665936261737 lags = 1.77071454279185e-07 wags = 1.23551824445621e-07 pags = -1.00320256456803e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.04518365194877+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.53043555901637e-07 wnfactor = -3.36356326968899e-07 pnfactor = 1.11774871374522e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.58153055902701 lpclm = -2.58735367075028e-06 wpclm = -6.73432761943568e-06 ppclm = 1.26598128421269e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 8.97336675484595e-06 lalpha0 = 1.03370180848787e-11 walpha0 = 3.78673832262507e-11 palpha0 = -7.12526315043093e-17   alpha1 = 0.0   beta0 = 23.755422300722 lbeta0 = 1.09371554517588e-05 wbeta0 = 3.6001833663671e-07 pbeta0 = -6.77423462875753e-13   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284635e-8   kt2 = -0.019151   at = 149419.117919288 lat = -0.269459747203754 wat = -0.0634618507974833 pat = 2.46335804682141e-7   ute = -1.22096728 lute = -1.46076520729919e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.36 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.765067508082857+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.62290355697613e-08 wvth0 = 5.0766518332166e-08 pvth0 = 9.29893193054649e-14   k1 = 0.88325   k2 = -0.0424095328288057 lk2 = 1.71927754471935e-08 wk2 = -4.40660856313329e-09 pk2 = -1.21272171837903e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 125882.1493544 lvsat = -0.0124492897266392 wvsat = -0.0819077852087622 pvsat = 9.42761751081294e-9   ua = -9.78864175812193e-10 lua = 7.33376932775916e-16 wua = 5.75680817817896e-15 pua = -5.09377167447714e-21   ub = 3.7197541520205e-18 lub = -1.38476205141157e-24 wub = -1.10966131451033e-23 pub = 9.18605229655207e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.038426162604325 lu0 = 7.01668748833791e-09 wu0 = 2.75549837343501e-08 pu0 = -3.12325498331512e-14   a0 = 1.56423106630244 la0 = 2.34069480918021e-08 wa0 = -2.12381543700583e-06 pa0 = -3.26805423624082e-13   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.230168630289976 lags = -5.53280301072259e-08 wags = -3.5675673647517e-07 pags = 8.03445622879953e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.894817092371182+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.01084242042997e-08 wnfactor = 1.73375496031912e-07 pnfactor = 1.58618965241267e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.142145193796235 lpclm = 1.21045650341096e-07 wpclm = -2.6859483867998e-06 ppclm = 5.04223673634689e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.91865203174779e-05 lalpha0 = -6.53294993320979e-11 walpha0 = -2.32289013861906e-10 palpha0 = 4.37083370887061e-16   alpha1 = 0.0   beta0 = 32.7578835350032 lbeta0 = -6.00219969526929e-06 wbeta0 = -4.16288555308075e-05 pbeta0 = 7.83303532055665e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 3474.80391928801 lat = 0.0051543280139506 wat = 0.0377190111718084 pat = 5.59502522896903e-8   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.1054288121068e-18 lub1 = -1.21755244170261e-24 wub1 = -4.46023452115792e-24 pub1 = 8.39253784345356e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.37 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.672532173788987+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.78115175552702e-08 wvth0 = 5.43325921797022e-07 pvth0 = -3.41268782927682e-13   k1 = 0.88325   k2 = -0.0192639554259554 lk2 = -3.21319883194586e-09 wk2 = -7.74231638401641e-08 pk2 = 5.22468065444297e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 169075.887664386 lvsat = -0.0505304443953024 wvsat = -0.581811391826307 pvsat = 4.50160633634678e-7   ua = -4.33199518312796e-09 lua = 3.68961794154176e-15 wua = 2.87693290946905e-14 pua = -2.53824385652267e-20   ub = 6.67586275993366e-18 lub = -3.9909738200577e-24 wub = -3.7542282609802e-23 pub = 3.25015065407312e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0194009801725477 lu0 = 2.37899732267604e-08 wu0 = 1.84649524927058e-07 pu0 = -1.69732752752126e-13   a0 = 3.1877872463121 la0 = -1.40797862822719e-06 wa0 = -1.09961878512208e-05 pa0 = 7.49539750215472e-12   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.191823757135535 lags = -2.15218095188377e-08 wags = 2.44458020380464e-06 pags = -1.66631387180058e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.768768221327417+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.10207982672393e-08 wnfactor = 6.5732606002195e-07 pnfactor = -2.68049274192641e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -3.94195754746114 lpclm = 3.72173765473228e-06 wpclm = 2.48882074952542e-05 ppclm = -1.92681317588837e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -0.000144860176257341 lalpha0 = 1.05749054049339e-10 walpha0 = 9.95115993328864e-10 palpha0 = -6.45041070032581e-16   alpha1 = 0.0   beta0 = -6.53739419501602 lbeta0 = 2.86419317815139e-05 wbeta0 = 0.000208144277654037 pbeta0 = -1.41878632842988e-10   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37954636 lkt1 = 6.00954836496102e-9   kt2 = -0.019151   at = -57748.01878932 lat = 0.059130572535477 wat = 0.446023452115794 pat = -3.04025641806401e-7   ute = -1.47412127 lute = 1.54745870397718e-7   ua1 = 6.387700286e-09 lua1 = -2.98283933094789e-15   ub1 = -1.32611871778042e-17 lub1 = 7.73612974079738e-24 wub1 = 1.13811572511505e-23 pub1 = -5.57380343311736e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.38 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.738872711960502+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.25914184781909e-08 wvth0 = 1.4540862551177e-07 pvth0 = -7.00340287569887e-14   k1 = 0.88325   k2 = -0.0189696305953616 lk2 = -3.41382123217239e-09 wk2 = -2.63804581462084e-09 pk2 = 1.27057783397074e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 54372.6150114965 lvsat = 0.0276554355627229 wvsat = 0.267885218778807 pvsat = -1.2902316523175e-7   ua = 3.87263145986975e-09 lua = -1.90295094488462e-15 wua = -2.88611407921912e-14 pua = 1.39005644065878e-20   ub = -3.56469055553775e-18 lub = 2.98935597968698e-24 wub = 3.45566759585809e-23 pub = -1.66437391819871e-29   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0715418649082754 lu0 = -1.17511308809622e-08 wu0 = -2.19344945894726e-07 pu0 = 1.05644422360952e-13   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.865427583899875+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.48657029992006e-08 wnfactor = 9.00039160282366e-07 pnfactor = -4.3349126100176e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.7029947195553 lpclm = -8.07701028747738e-07 wpclm = -1.15171677732429e-05 ppclm = 5.54708261763362e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -7.46866227004865e-06 lalpha0 = 1.20980520210972e-11 walpha0 = 1.66329075980662e-10 palpha0 = -8.01100708390223e-17   alpha1 = 0.0   beta0 = 31.92270996 lbeta0 = 2.42614022570543e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10799999995 lat = 0.015430120515312   ute = -1.12187464 lute = -8.535811348896e-8   ua1 = 2.0117e-9   ub1 = -3.2720457516618e-18 lub1 = 9.27171335647382e-25 wub1 = 1.09200153546392e-23 pub1 = -5.25947251534701e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.39 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.760960415803883+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.19531851498796e-08 wvth0 = -1.29357769119043e-08 pvth0 = 6.23033584874137e-15   k1 = 0.88325   k2 = 0.0140043162181216 lk2 = -1.92952610796312e-08 wk2 = -1.72108259314386e-07 pk2 = 8.28935335831437e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 119417.903431542 lvsat = -0.003672716970754 wvsat = -0.0867469338286195 pvsat = 4.17804462214811e-8   ua = 1.95734028973037e-10 lua = -1.32024773857258e-16 wua = -2.59005145183813e-17 pua = 1.2474620210576e-23   ub = -1.14271444709589e-18 lub = 1.82284509472147e-24 wub = 2.96686226685909e-24 pub = -1.42894767476092e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0279896066426879 lu0 = 9.22520458104242e-09 wu0 = 2.21967634672392e-08 pu0 = -1.06907603693068e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {-0.289171459834467+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.31230762028834e-07 wnfactor = 5.6318897391071e-06 pnfactor = -2.71252084638458e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.0383260320000041 lpclm = 4.75699339251646e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.979747388e-05 lalpha0 = -5.85066072966767e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.447057200000001 lkt1 = 3.67619272991999e-8   kt2 = -0.019151   at = 121925.612125824 lat = -0.0402289417218334 wat = -0.617828151016205 pat = 2.97568279342841e-7   ute = -1.30100818 lute = 9.19048182478768e-10   ua1 = -1.77680057200001e-09 lua1 = 1.82467826149579e-15   ub1 = 7.06998198e-18 lub1 = -4.05392153291928e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.40 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.786974616656+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.37021580860907e-8   k1 = 0.88325   k2 = -0.042883449483 wk2 = 1.04535575894407e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 132252.653514 wvsat = -0.156881217012554   ua = 3.825241555083e-10 wua = -1.53432816969018e-15   ub = 1.11223625989e-18 wub = 2.00358674204115e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04501150807589 wu0 = -1.28876015911906e-8   a0 = 0.6274899071701 wa0 = 9.60128477199801e-7   keta = -0.012522079359 wketa = -5.15175664817461e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.115611889898 wags = 1.70838167294462e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.03539243781+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -6.64582977419424e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.79888786264 wpclm = 4.91295974020729e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.265792481e-06 walpha0 = 2.66187069017512e-11   alpha1 = 0.0   beta0 = 21.634866085 wbeta0 = 6.26364148047058e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 207544.7936 wat = -0.271778342203469   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.41 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.786974616656+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.37021580860924e-8   k1 = 0.88325   k2 = -0.042883449483 wk2 = 1.04535575894406e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 132252.653514 wvsat = -0.156881217012554   ua = 3.825241555083e-10 wua = -1.53432816969018e-15   ub = 1.11223625989e-18 wub = 2.00358674204114e-24   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.04501150807589 wu0 = -1.28876015911906e-8   a0 = 0.6274899071701 wa0 = 9.601284771998e-7   keta = -0.012522079359 wketa = -5.15175664817461e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.115611889898 wags = 1.70838167294462e-7   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.03539243781+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -6.64582977419407e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.79888786264 wpclm = 4.91295974020729e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.265792481e-06 walpha0 = 2.66187069017512e-11   alpha1 = 0.0   beta0 = 21.634866085 wbeta0 = 6.26364148047058e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.40273   kt2 = -0.019151   at = 207544.7936 wat = -0.271778342203469   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.42 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.786357685474902+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.86242700646278e-09 wvth0 = 3.08403082604422e-09 pvth0 = 8.3688214065364e-14   k1 = 0.88325   k2 = -0.0419646716003985 lk2 = -7.24147283551573e-09 wk2 = 4.39586791068118e-09 pk2 = 4.77445050489397e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 137283.136891999 lvsat = -0.0396484388894403 wvsat = -0.193982849262734 pvsat = 2.92421560401781e-7   ua = 3.84047811182946e-10 lua = -1.20088994168929e-17 wua = -1.54004932105345e-15 pua = 4.50920325462213e-23   ub = 9.46525747431211e-19 lub = 1.30606994057364e-24 wub = 2.00441091750764e-24 pub = -6.49585102706769e-33   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0433619005933727 lu0 = 1.30016057200779e-08 wu0 = -9.96363307992266e-09 pu0 = -2.30456554812755e-14   a0 = 0.634468848653946 la0 = -5.50054764409682e-08 wa0 = 9.54662133418256e-07 pa0 = 4.30837319370173e-14   keta = -0.012522079359 wketa = -5.15175664817461e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.104497467101648 lags = 8.75998348309459e-08 wags = 1.22095056579999e-07 pags = 3.84175456159097e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.12202402115767+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.82798606050028e-07 wnfactor = -1.22502229463798e-07 pnfactor = 4.4171786984053e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.798887862639999 wpclm = 4.91295974020729e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -7.22268727179076e-06 lalpha0 = 9.84296516048668e-11 walpha0 = 6.43728113962422e-11 palpha0 = -2.97564109131542e-16   alpha1 = 0.0   beta0 = 16.9309081340308 lbeta0 = 3.70748843288447e-05 wbeta0 = 1.17306720749066e-05 pbeta0 = -4.30891451462084e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.414374908 lkt1 = 9.17809261094877e-8   kt2 = -0.019151   at = 303241.884414362 lat = -0.754249636057748 wat = -0.398151913733146 pat = 9.96030490816877e-7   ute = -1.33741636 lute = 3.05936420364961e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.43 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.793270887647352+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.19721074213994e-08 wvth0 = -1.00544015368319e-08 pvth0 = 1.34686826108684e-13   k1 = 0.88325   k2 = -0.0490118449921127 lk2 = 2.0113089100004e-08 wk2 = 1.93647720563838e-08 pk2 = -1.03593321635693e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 144500.64632635 lvsat = -0.0676641833401563 wvsat = -0.207302121448226 pvsat = 3.44122126810781e-7   ua = 4.57074803764835e-10 lua = -2.95473102794488e-16 wua = -1.74251532275337e-15 pua = 8.30991353520685e-22   ub = 1.17391334069664e-18 lub = 4.23434072601203e-25 wub = 2.43804973671967e-24 pub = -1.68972390267799e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0462217969917336 lu0 = 1.90052890392952e-09 wu0 = -1.77986599767687e-08 pu0 = 7.36706698249045e-15   a0 = 0.166730231382506 la0 = 1.76058557895007e-06 wa0 = 1.85263333213487e-06 pa0 = -3.44251359996455e-12   keta = -0.0410423384854744 lketa = 1.10705264554652e-07 wketa = 3.09903453202611e-08 pketa = -3.20265680735496e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.0357471351464282 lags = 3.54463598360278e-07 wags = 4.70522375147385e-07 pags = -9.68292566975537e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.01837925571955+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.80487353313839e-07 wnfactor = -2.05203542003951e-07 pnfactor = 7.62734261843633e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.798887862640001 wpclm = 4.91295974020729e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.1586090330971e-05 lalpha0 = -1.33955366540069e-11 walpha0 = -2.38461434973391e-11 palpha0 = 4.48697620657591e-17   alpha1 = 0.0   beta0 = 24.0309567985967 lbeta0 = 9.51507983071382e-06 wbeta0 = -9.88160389015598e-07 pbeta0 = 6.28073282372086e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.5734434328464e-8   kt2 = -0.019151   at = 178987.39479822 lat = -0.271938936002104 wat = -0.208138187698469 pat = 2.58466371346539e-7   ute = -1.22096728 lute = -1.46076520729921e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.44 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.759391035323052+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.17774423866912e-08 wvth0 = 7.85412611340402e-08 pvth0 = -3.20179622166859e-14   k1 = 0.88325   k2 = -0.0476279347631974 lk2 = 1.75090737925088e-08 wk2 = 2.1126812928964e-08 pk2 = -1.36748517028874e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123496.862325666 lvsat = -0.0281427072282449 wvsat = -0.0702366759592215 pvsat = 8.62148502226343e-8   ua = 7.01032121160565e-10 lua = -7.54511973669719e-16 wua = -2.46285384726428e-15 pua = 2.18640625342729e-21   ub = 7.78802199614433e-19 lub = 1.16688941966257e-24 wub = 3.29334123803762e-24 pub = -3.29907118205187e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.047592351445367 lu0 = -6.78355695987298e-10 wu0 = -1.72947932849368e-08 pu0 = 6.41897327593861e-15   a0 = 1.12961416130036 la0 = -5.12114874048397e-08 wa0 = 2.74682525933684e-09 pa0 = 3.82994472867002e-14   keta = 0.0428767626961974 lketa = -4.71999373164247e-08 wketa = -2.61953131328461e-07 pketa = 2.30947310891899e-13   a1 = 0.0   a2 = 0.65972622   ags = 0.156710711342347 lags = 1.26854178701294e-07 wags = 2.66977570298117e-09 pags = -8.79642731673668e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.862589222006669+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.26527825615269e-08 wnfactor = 3.31065112154916e-07 pnfactor = -2.4632814349324e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.29612431526648 lpclm = 2.81725400977428e-06 wpclm = 9.24440191372468e-06 ppclm = -8.15019752560857e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.12022666393148e-05 lalpha0 = 4.83002162021337e-11 walpha0 = 6.31907843886289e-11 palpha0 = -1.18902054773882e-16   alpha1 = 0.0   beta0 = 21.3097487258468 lbeta0 = 1.46354029038908e-05 wbeta0 = 1.43863872687332e-05 pbeta0 = -2.26485695328151e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 30749.501838576 lat = 0.00699081995490923 wat = -0.0957349402099551 pat = 4.69643743552413e-8   ute = -1.2986   ua1 = 3.0044e-9   ub1 = -4.0169908e-18 lub1 = 4.97675410948802e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.45 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.745533355563818+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.39948717389003e-08 wvth0 = 1.86134205422418e-07 pvth0 = -1.26875775247315e-13   k1 = 0.88325   k2 = -0.0401469672038876 lk2 = 1.09135834773891e-08 wk2 = 2.47565357027634e-08 pk2 = -1.68749459702888e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 25344.8904415296 lvsat = 0.0583916046557976 wvsat = 0.121458340883249 pvsat = -8.27903776462942e-8   ua = 1.53235127150898e-09 lua = -1.4874328641063e-15 wua = 7.53281947029906e-17 pua = -5.1346409324568e-23   ub = -5.92658179390834e-19 lub = 2.37601826236725e-24 wub = -1.97771493156669e-24 pub = 1.34808169509339e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0661606744945015 lu0 = -1.70488577557341e-08 wu0 = -4.41436954831001e-08 pu0 = 3.00899320143184e-14   a0 = 0.898825520536816 la0 = 1.52260086683369e-07 wa0 = 2.03605736605214e-07 pa0 = -1.38784999876633e-13   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.778919072031579 lags = -4.21707111583317e-07 wags = -4.28052513978468e-07 pags = 2.91776003418227e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.856562183872992+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.79664363535485e-08 wnfactor = 2.27753888632863e-07 pnfactor = -1.55245249632146e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.144578551 lpclm = -2.16193502429436e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 0.000123090195536574 lalpha0 = -7.00968529807682e-11 walpha0 = -3.15953921943145e-10 palpha0 = 2.15365567537637e-16   alpha1 = 0.0   beta0 = 46.1851798977574 lbeta0 = -7.29567273278776e-06 wbeta0 = -4.98250630337912e-05 pbeta0 = 3.39625566661012e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.379546360000001 lkt1 = 6.00954836496017e-9   kt2 = -0.019151   at = 71666.21878932 lat = -0.0290828307106769 wat = -0.187194976958514 pat = 1.27598835314093e-7   ute = -1.47412127 lute = 1.54745870397719e-7   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -1.093515919e-17 lub1 = 6.59698171763484e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.46 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.81191695338626+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.74542165360274e-09 wvth0 = -2.11993779926313e-07 pvth0 = 1.44502592173854e-13   k1 = 0.88325   k2 = -0.0130220285453547 lk2 = -7.5757512100586e-09 wk2 = -3.17394128460188e-08 pk2 = 2.16347264147089e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 106894.824168398 lvsat = 0.00280423402994989 wvsat = 0.0108962553068732 pvsat = -7.42727988235601e-9   ua = -2.2598777560032e-09 lua = 1.097486961291e-15 wua = 1.14496923568805e-15 pua = -7.80452249937461e-22   ub = 2.97916661184504e-18 lub = -5.86661010316081e-26 wub = 2.53785768057792e-24 pub = -1.72989515795841e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0205531526180277 lu0 = 1.4038871026058e-08 wu0 = 3.01406818155405e-08 pu0 = -2.05449737900177e-14   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.12147940482315+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.62610678466036e-07 wnfactor = -3.52811645318757e-07 pnfactor = 2.40489118668497e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.25066874317934 lpclm = -2.88508396665789e-07 wpclm = -4.4109977685263e-06 ppclm = 3.00669487494719e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.85382953993712e-05 lalpha0 = -5.64687397884577e-12 walpha0 = -9.85145560358655e-12 palpha0 = 6.71510679180632e-18   alpha1 = 0.0   beta0 = 31.92270996 lbeta0 = 2.42614022570543e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000004 lat = 0.015430120515312   ute = -1.12187464 lute = -8.53581134889591e-8   ua1 = 2.0117e-9   ub1 = -1.61850517850452e-18 lub1 = 2.46414943855107e-25 wub1 = 2.82931077888471e-24 pub1 = -1.92856008207586e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.47 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.760165258917606+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.36709007707086e-08 wvth0 = -9.0451076639278e-09 pvth0 = 4.67552054600853e-14   k1 = 0.88325   k2 = -0.0506406950412919 lk2 = 1.05427528463786e-08 wk2 = 1.44197065687451e-07 pk2 = -6.31026153602376e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 128991.278447869 lvsat = -0.00783821382339739 wvsat = -0.133589055701759 pvsat = 6.2162047370598e-8   ua = 6.70040009111595e-10 lua = -3.13666911427831e-16 wua = -2.34665975448518e-15 pua = 9.01241970373615e-22   ub = -8.69696500986132e-19 lub = 1.79508493317995e-24 wub = 1.63099692329779e-24 pub = -1.29311837026504e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0330807201115519 lu0 = 8.00514352874704e-09 wu0 = -2.713840909148e-09 pu0 = -4.7210528829897e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.674356934717602+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.27395995457223e-08 wnfactor = 9.17385772756392e-07 pnfactor = -3.71283684983545e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.76467238675867 lpclm = 1.16378844379303e-06 wpclm = 8.82199553705259e-06 ppclm = -3.3667910887786e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.57706845212577e-05 lalpha0 = -4.3138929459547e-12 walpha0 = 1.97029112071731e-11 palpha0 = -7.51934022146076e-18   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4470572 lkt1 = 3.67619272991999e-8   kt2 = -0.019151   at = -4343.23199999996 lat = 0.020586679287552   ute = -1.30100818 lute = 9.19048182479615e-10   ua1 = -1.776800572e-09 lua1 = 1.82467826149579e-15   ub1 = 8.22646473700904e-18 lub1 = -4.49527698637318e-24 wub1 = -5.65862155776943e-24 pub1 = 2.1595336968209e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.48 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.780586837412+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.21817351522552e-8   k1 = 0.88325   k2 = -0.0420744887733333 wk2 = 8.11326823272488e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 42590.8630346667 wvsat = 0.102506577048957   ua = -1.48366523663467e-10 wua = 1.5162677452152e-18   ub = 1.66245897878667e-18 wub = 4.11815525627282e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0412881053152787 wu0 = -2.11595378765795e-9   a0 = 0.8146724514104 wa0 = 4.18617238379473e-7   keta = -0.0348366834493333 wketa = 1.30376459382165e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.155519256609333 wags = 5.53878315079763e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.07611532614667+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.84267903338609e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.32650592750667 wpclm = -1.23571522814783e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.1069478666667 wbeta0 = 7.79088671354373e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.413873664 wkt1 = 3.22381519181116e-8   kt2 = -0.019151   at = 154088.645866667 wat = -0.11713195196914   ute = -1.405857766 wute = 3.10292212211828e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.49 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.780586837412+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.21817351522548e-8   k1 = 0.88325   k2 = -0.0420744887733333 wk2 = 8.11326823272485e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 42590.8630346666 wvsat = 0.102506577048957   ua = -1.48366523663467e-10 wua = 1.5162677452152e-18   ub = 1.66245897878667e-18 wub = 4.11815525627282e-25   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0412881053152787 wu0 = -2.11595378765795e-9   a0 = 0.8146724514104 wa0 = 4.18617238379473e-7   keta = -0.0348366834493333 wketa = 1.30376459382165e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.155519256609333 wags = 5.53878315079763e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.07611532614667+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.84267903338609e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.32650592750667 wpclm = -1.23571522814783e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.4467e-5   alpha1 = 0.0   beta0 = 21.1069478666667 wbeta0 = 7.79088671354373e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.413873664 wkt1 = 3.22381519181116e-8   kt2 = -0.019151   at = 154088.645866667 wat = -0.11713195196914   ute = -1.405857766 wute = 3.10292212211828e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.50 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.772318248574765+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.51700074487538e-08 wvth0 = 4.36995321217929e-08 pvth0 = -9.07790832358024e-14   k1 = 0.88325   k2 = -0.0443409580087096 lk2 = 1.78634855184343e-08 wk2 = 1.12703646858961e-08 pk2 = -2.48830850607871e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 27558.4262893798 lvsat = 0.118480194619376 wvsat = 0.123446130072798 pvsat = -1.65037934936616e-7   ua = -1.49242043323507e-10 lua = 6.90052727128287e-18 wua = 2.73582985982581e-18 pua = -9.61214466675168e-24   ub = 1.3434127272965e-18 lub = 2.51460642140998e-24 wub = 8.56233554010527e-25 pub = -3.50274113155441e-30   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0400559208805184 lu0 = 9.71162919964623e-09 wu0 = -3.99572621783156e-10 pu0 = -1.35278915866807e-14   a0 = 0.824488078620849 la0 = -7.73632007844582e-08 wa0 = 4.04944481931658e-07 pa0 = 1.07763689438317e-13   keta = -0.0348366834493333 wketa = 1.30376459382165e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.101588143903633 lags = 4.25065399421306e-07 wags = 1.30511606400284e-07 pags = -5.92098248647105e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.20583372639764+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.0223932132805e-06 wnfactor = -3.64960186715407e-07 pnfactor = 1.42415080558477e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.32650592750667 wpclm = -1.23571522814783e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.55506380572113e-05 lalpha0 = -8.54084072268658e-12 walpha0 = -1.50946230089693e-12 palpha0 = 1.18970324113921e-17   alpha1 = 0.0   beta0 = 15.6793997390108 lbeta0 = 4.27779587146651e-05 wbeta0 = 1.5351233298347e-05 pbeta0 = -5.95878998152624e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.436332483838576 lkt1 = 1.77012242957235e-07 wkt1 = 6.35223446828149e-08 pkt1 = -2.46570619925222e-13   kt2 = -0.019151   at = 254404.707812306 lat = -0.790654685208982 wat = -0.256868012984814 pat = 1.10134876899933e-6   ute = -1.48072049879525 lute = 5.90040809857453e-07 wute = 4.14572854760838e-07 pute = -8.21902066417413e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.51 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.782053190287529+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.73825072385864e-08 wvth0 = 2.2397925781847e-08 pvth0 = -8.09400120883733e-15   k1 = 0.88325   k2 = -0.0444199778610054 lk2 = 1.81702118218201e-08 wk2 = 6.08069330451002e-09 pk2 = -4.73866979862897e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 28186.7954070382 lvsat = 0.116041094430984 wvsat = 0.129188964079605 pvsat = -1.87329526159462e-7   ua = -1.4499904126515e-10 lua = -9.56926226651178e-18 wua = -7.4097618311703e-19 pua = 3.8835508345534e-24   ub = 2.05010293237498e-18 lub = -2.2850771947006e-25 wub = -9.67299520429297e-26 pub = 1.96316320228907e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0414400102869553 lu0 = 4.33909793240191e-09 wu0 = -3.96515187488666e-09 pu0 = 3.12389203018964e-16   a0 = 0.516408528979551 la0 = 1.11848946996699e-06 wa0 = 8.4102870367512e-07 pa0 = -1.58495652471308e-12   keta = -0.0272933305616225 lketa = -2.92805501296425e-08 wketa = -8.78495714510981e-09 pketa = 8.47074017419502e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.21163507679463 lags = -2.09673697797468e-09 wags = -3.8314052747315e-08 pags = 6.3221507623943e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.951889578982612+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.66744686850067e-08 wnfactor = -1.28516997704185e-08 pnfactor = 5.73938267535807e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.32650592750667 wpclm = -1.23571522814783e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.12888761567053e-05 lalpha0 = 8.00176769374573e-12 walpha0 = 5.94326462581616e-12 palpha0 = -1.70317407255068e-17   alpha1 = 0.0   beta0 = 22.7536711488142 lbeta0 = 1.53182121366015e-05 wbeta0 = 2.70697334980803e-06 pbeta0 = -1.05074852056554e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.5734434328464e-8   kt2 = -0.019151   at = 97754.5133333333 lat = -0.1825956509124 wat = 0.0268651265984267 pat = 1.05879118406788e-22   ute = -1.26626698809741 lute = -2.42389657593698e-07 wute = 1.31050152938058e-07 pute = 2.78629859795158e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.52 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.782622293562378+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.63116620289116e-08 wvth0 = 1.13342067605102e-08 pvth0 = 1.27238907955936e-14   k1 = 0.88325   k2 = -0.0408057828744032 lk2 = 1.136961242401e-08 wk2 = 1.39061404506183e-09 pk2 = 4.08635217880209e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 81623.3624165292 lvsat = 0.015492926229514 wvsat = 0.0509016005909145 pvsat = -4.00212046740568e-8   ua = -1.5057461334727e-10 lua = 9.21934883800956e-19 wua = 8.0866818404126e-19 pua = 9.67684206111081e-25   ub = 1.86521434079331e-18 lub = 1.19385310439315e-25 wub = 1.50396542917043e-25 pub = -2.68685789241595e-31   uc = 6.6204e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0428247204684782 lu0 = 1.73357740528203e-09 wu0 = -3.50223710929852e-09 pu0 = -5.58647884843313e-16   a0 = 1.13446565679043 la0 = -4.44690717785511e-08 wa0 = -1.12883474306116e-08 pa0 = 1.87939220613015e-14   keta = -0.0712384237142915 lketa = 5.34081191697731e-08 wketa = 6.81773101192543e-08 pketa = -6.01075709842989e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.150292596396241 lags = 1.1332748246893e-07 wags = 2.12371126812386e-08 pags = -4.88321090883785e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.977525230672974+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.49114337890532e-08 wnfactor = -1.4399336043415e-09 pnfactor = 3.5921036711904e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.91345540001117 lpclm = -1.10442525764549e-06 wpclm = -2.93373540022552e-06 ppclm = 3.19505588450758e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.00063250950864e-05 lalpha0 = -8.4012980568738e-12 walpha0 = -2.70943607381408e-11 palpha0 = 4.51330445138278e-17   alpha1 = 0.0   beta0 = 29.3649587667896 lbeta0 = 2.87817534826473e-06 wbeta0 = -8.91699706089276e-06 pbeta0 = 1.1364595982054e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = -19816.50346192 lat = 0.0386302068461533 wat = 0.0505503893521571 pat = -4.45670430668784e-8   ute = -1.48015069840935 lute = 1.60061631542824e-07 wute = 5.25218545368912e-07 pute = -4.63051577464866e-13   ua1 = 3.0044e-9   ub1 = -4.2626071838576e-18 lub1 = 9.59836041005078e-25 wub1 = 7.10557882611913e-25 pub1 = -1.33701129200635e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.53 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.845770510427469+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.93620792951599e-08 wvth0 = -1.0384767363762e-07 pvth0 = 1.1427238310228e-13   k1 = 0.88325   k2 = -0.0258848913074395 lk2 = -1.78518273352157e-09 wk2 = -1.6503050858473e-08 pk2 = 1.98620513296949e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93101.377072713 lvsat = 0.00537349530009457 wvsat = -0.0745583291683265 pvsat = 7.05887859591615e-8   ua = 3.16755375719576e-09 lua = -2.92445948920827e-15 wua = -4.65524391788445e-15 pua = 4.10591126197719e-21   ub = -3.99386674728161e-18 lub = 5.28496212460534e-24 wub = 7.86183860458147e-24 pub = -7.06737072271917e-30   uc = 6.49475078108089e-11 luc = 1.10776874770968e-18 wuc = 3.63497913065784e-18 puc = -3.20472846083672e-24   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0558722625567314 lu0 = -9.76960541123715e-09 wu0 = -1.43797518604327e-08 pu0 = 9.0313607102876e-15   a0 = 0.953923864057659 la0 = 1.14703072199193e-07 wa0 = 4.42085429298374e-08 pa0 = -3.01341343685228e-14   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.68299338492663 lags = -3.56320709927849e-07 wags = -1.50543530062711e-07 pags = 1.02615889657826e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.0533658523146+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.51775256090693e-07 wnfactor = -3.41590858414642e-07 pnfactor = 3.35810337457959e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.726995206800878 lpclm = -5.83992387443388e-08 wpclm = 1.2080510762676e-06 ppclm = -4.56492177481913e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.56417217617624e-05 lalpha0 = -4.55330663249543e-12 walpha0 = -5.11000014851337e-12 palpha0 = 2.57508407810309e-17   alpha1 = 0.0   beta0 = 27.585680224269 lbeta0 = 4.44685136537833e-06 wbeta0 = 3.98250834262432e-06 pbeta0 = -8.07236388120435e-15   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37954636 lkt1 = 6.00954836495975e-9   kt2 = -0.019151   at = 6959.10000000001 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397719e-7   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -1.14294527099004e-17 lub1 = 7.27838506320338e-24 wub1 = 1.42997039274411e-24 pub1 = -1.97127125978927e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.54 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.720733715736931+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.58675012905208e-08 wvth0 = 5.17954968972161e-08 pvth0 = 8.18039491159715e-15   k1 = 0.88325   k2 = -0.0296782071230875 lk2 = 8.00477885793404e-10 wk2 = 1.64462122198618e-08 pk2 = -2.59735255796894e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 94534.8384209295 lvsat = 0.00439639644054179 wvsat = 0.0466531749548986 pvsat = -1.20333388653772e-8   ua = -3.46057585700204e-09 lua = 1.59351226849506e-15 wua = 4.61853841255745e-15 pua = -2.2154326306159e-21   ub = 7.2786586550529e-18 lub = -2.39879700054035e-24 wub = -9.9003922217566e-24 pub = 5.0400052488226e-30   uc = 5.20633665815315e-11 luc = 9.89006323866942e-18 wuc = 4.09082585730258e-17 puc = -2.86115375668146e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0307387566130352 lu0 = 7.36229704620009e-09 wu0 = 6.74157253351747e-10 pu0 = -1.22992568239593e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.832672495537658+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.34271915068245e-09 wnfactor = 4.82694613353996e-07 pnfactor = -2.26052314376529e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.126006858428593 lpclm = 3.51256055086753e-07 wpclm = -1.15739817174156e-06 ppclm = 1.15588318613406e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.01170667724411e-05 lalpha0 = 1.3004810948805e-11 walpha0 = 1.01976883634255e-10 palpha0 = -4.72434343331203e-17   alpha1 = 0.0   beta0 = 27.2448876536411 lbeta0 = 4.67914785005091e-06 wbeta0 = 1.35327434637594e-05 pbeta0 = -6.51785643091123e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000004 lat = 0.015430120515312   ute = -1.12187464 lute = -8.535811348896e-8   ua1 = 2.0117e-9   ub1 = 4.37359482859094e-19 lub1 = -8.10461332620454e-25 wub1 = -3.11821934012444e-24 pub1 = 1.12893859696432e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.55 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.737449143880527+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.78167493411504e-08 wvth0 = 5.66716590615061e-08 pvth0 = 5.83185967143656e-15   k1 = 0.88325   k2 = -0.0163946867859807 lk2 = -5.59734371528934e-09 wk2 = 4.51248021371831e-08 pk2 = -1.64099938913879e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 71665.6049018061 lvsat = 0.0154110425957582 wvsat = 0.0322517101887114 pvsat = -5.09707498124991e-9   ua = -1.67314729107859e-10 lua = 7.35915190061682e-18 wua = 7.57723342846933e-17 pua = -2.74729477409262e-23   ub = -2.64449019184359e-18 lub = 2.38054871748349e-24 wub = 6.76540052961341e-24 pub = -2.98684050877625e-30   uc = 9.6998251215319e-11 luc = -1.17521948568096e-17 wuc = -8.90864754073672e-17 puc = 3.3998606128566e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0268075249178557 lu0 = 9.25571975493955e-09 wu0 = 1.54342493120171e-08 pu0 = -8.33891738116328e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.20891981211057+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.82556971715595e-07 wnfactor = -6.29082179900626e-07 pnfactor = 3.09419413219455e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.783804384471329 lpclm = 7.89453902872101e-07 wpclm = 5.98438560289141e-06 ppclm = -2.28385698394507e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.61093936479351e-05 lalpha0 = -4.44315654222335e-12 walpha0 = 1.87230399294786e-11 palpha0 = -7.14538606652652e-18   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4470572 lkt1 = 3.67619272992001e-8   kt2 = -0.019151   at = -4343.23200000008 lat = 0.020586679287552   ute = -1.30100818 lute = 9.19048182480462e-10   ua1 = -1.776800572e-09 lua1 = 1.82467826149579e-15   ub1 = 6.85068240027468e-18 lub1 = -3.89934852927283e-24 wub1 = -1.67854104045507e-24 pub1 = 4.35537699424768e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.56 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.800086021512+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.02019066668706e-9   k1 = 0.88325   k2 = -0.037600152496 wk2 = 1.88070572052318e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123823.72048 wvsat = -0.0106473815923799   ua = -1.47610180376e-10 wua = 4.62713312192173e-19   ub = 2.22289776532e-18 wub = -3.68852165584617e-25   uc = 9.0417449128e-11 wuc = -3.37283176704406e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.042547130988724 wu0 = -3.869723671689e-9   a0 = 1.1095237950092 wa0 = 7.90170050277481e-9   keta = -0.031975948324 wketa = 9.05276205950239e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.2281875023 wags = -4.58359826728035e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.80418922796+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.94513730539294e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.611460833560001 wpclm = 1.46379107541407e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.4729154768e-05 walpha0 = 4.06690173533238e-11   alpha1 = 0.0   beta0 = 26.224946344 wbeta0 = 6.61729790554457e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.387158168 wkt1 = -4.97541195905582e-9   kt2 = -0.019151   at = -72873.2800000001 wat = 0.19901647836224   ute = -1.2088171904 wute = 3.58229661052034e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.57 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.800086021512+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.02019066668706e-9   k1 = 0.88325   k2 = -0.037600152496 wk2 = 1.88070572052318e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123823.72048 wvsat = -0.0106473815923798   ua = -1.47610180376e-10 wua = 4.62713312192271e-19   ub = 2.22289776532e-18 wub = -3.68852165584616e-25   uc = 9.0417449128e-11 wuc = -3.37283176704407e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.042547130988724 wu0 = -3.869723671689e-9   a0 = 1.1095237950092 wa0 = 7.90170050277524e-9   keta = -0.031975948324 wketa = 9.0527620595024e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.2281875023 wags = -4.58359826728035e-8   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.804189227959999+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.94513730539294e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.611460833560002 wpclm = 1.46379107541407e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -1.4729154768e-05 walpha0 = 4.06690173533238e-11   alpha1 = 0.0   beta0 = 26.224946344 wbeta0 = 6.61729790554457e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.387158168 wkt1 = -4.97541195905603e-9   kt2 = -0.019151   at = -72873.2800000001 wat = 0.19901647836224   ute = -1.2088171904 wute = 3.58229661052026e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.58 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.812394277263393+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.70091916273779e-08 wvth0 = -1.21246926482594e-08 pvth0 = 1.35129729550887e-13   k1 = 0.88325   k2 = -0.0340052475530105 lk2 = -2.83337322152444e-08 wk2 = -3.12684587905367e-09 pk2 = 3.94676989590824e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123823.72048 wvsat = -0.0106473815923798   ua = -1.4068795633739e-10 lua = -5.45584501827745e-17 wua = -9.17965404018204e-18 pua = 7.5997629649697e-23   ub = 3.15951755387e-18 lub = -7.3820962437481e-24 wub = -1.67352419300365e-24 pub = 1.02829500194989e-29   uc = 9.04174491280001e-11 wuc = -3.37283176704407e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0451351228661604 lu0 = -2.03976099489101e-08 wu0 = -7.47468766129901e-09 pu0 = 2.84130139592139e-14   a0 = 1.09286778915875 la0 = 1.3127657532712e-07 wa0 = 3.11028171002065e-08 pa0 = -1.82862755814517e-13   keta = -0.031975948324 wketa = 9.0527620595024e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.322365935704974 lags = -7.42280131148247e-07 wags = -1.77022584911729e-07 pags = 1.033965046924e-12   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.767188205671601+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.91628589305052e-07 wnfactor = 2.46054600544098e-07 pnfactor = -4.06226376501183e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.611460833560001 wpclm = 1.46379107541407e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -3.05243452661954e-05 lalpha0 = 1.24491942057435e-10 walpha0 = 6.26710543193091e-11 palpha0 = -1.7341204662444e-16   alpha1 = 0.0   beta0 = 28.1729158546399 lbeta0 = -1.53531866219614e-05 wbeta0 = -2.05170992304739e-06 pbeta0 = 2.13863441305541e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.383692030080713 lkt1 = -2.73188374056248e-08 wkt1 = -9.8035965028316e-09 pkt1 = 3.80539931148653e-14   kt2 = -0.019151   at = -263510.86556084 lat = 1.5025360573094 wat = 0.464566628269897 pat = -2.09296962131758e-6   ute = -1.2088171904 wute = 3.58229661052026e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.59 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.773909346029202+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.23753029087767e-08 wvth0 = 3.37419587922368e-08 pvth0 = -4.29079158799944e-14   k1 = 0.88325   k2 = -0.0451283325544879 lk2 = 1.48420349575507e-08 wk2 = 7.06740164163409e-09 pk2 = -1.0265921013003e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 133867.550425757 lvsat = -0.0389864918953293 wvsat = -0.0180198890697598 pvsat = 2.86173904344667e-8   ua = -1.53450450871192e-10 lua = -5.0190919505639e-18 wua = 1.1031482438897e-17 pua = -2.45464530840874e-24   ub = 5.10719696666901e-19 lub = 2.89957287549432e-24 wub = 2.04756624120253e-24 pub = -4.16096856917148e-30   uc = 1.12530849807749e-10 luc = -8.58361721609397e-17 wuc = -6.4531356054503e-17 puc = 1.19566182700958e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0371451450807145 lu0 = 1.06165754622768e-08 wu0 = 2.0174149730682e-09 pu0 = -8.43187334204058e-15   a0 = 1.14498129709505 la0 = -7.1009093164701e-08 wa0 = -3.45467622535062e-08 pa0 = 7.19650147897095e-14   keta = -0.0546060069871326 lketa = 8.78416503889275e-08 wketa = 2.9260453983216e-08 pketa = -7.84389044479959e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.0539739199129321 lags = 2.99519979462711e-07 wags = 1.81301317020302e-07 pags = -3.56917910475841e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.745564095251705+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.75565514778891e-07 wnfactor = 2.74551033396416e-07 pnfactor = -5.16839156132324e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.611460833560002 wpclm = 1.46379107541407e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -6.60165003024548e-06 lalpha0 = 3.1632747012543e-11 walpha0 = 3.08640162021387e-11 palpha0 = -4.994870241546e-17   alpha1 = 0.0   beta0 = 21.1207507685435 lbeta0 = 1.20207512541732e-05 wbeta0 = 4.98156285686912e-06 pbeta0 = -5.91426068978983e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284635e-8   kt2 = -0.019151   at = 221025.03757864 lat = -0.378255947609322 wat = -0.144845536313267 pat = 2.72546575566351e-7   ute = -1.17841312733626 lute = -1.18017505734487e-07 wute = 8.67341475993078e-09 pute = 1.05384675885656e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.60 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.78370312202232+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.39469814241918e-08 wvth0 = 9.82865811060713e-09 pvth0 = 2.08821156138247e-15   k1 = 0.88325   k2 = -0.0484860500256003 lk2 = 2.11600370290247e-08 wk2 = 1.2088903615459e-08 pk2 = -9.55129809815e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 128969.405699254 lvsat = -0.0297699664447308 wvsat = -0.0150494491681034 pvsat = 2.30281037796738e-8   ua = -1.63961328849154e-10 lua = 1.4758554444376e-17 wua = 1.94558006361142e-17 pua = -1.83061457037483e-23   ub = 2.097976425773e-18 lub = -8.70665272339636e-26 wub = -1.73831265452094e-25 pub = 1.88929496600975e-32   uc = 3.62663988019567e-11 luc = 5.76657643717961e-17 wuc = 4.1701821089624e-17 puc = -8.03259878078083e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0431773458390532 lu0 = -7.338306438406e-10 wu0 = -3.99342944024394e-09 pu0 = 2.87834789644645e-15   a0 = 1.1027916786562 la0 = 8.37641171611032e-09 wa0 = 3.28321738032901e-08 pa0 = -5.48176169364534e-14   keta = -0.00550873841431287 lketa = -4.54153765935886e-09 wketa = -2.33813808568333e-08 pketa = 2.06138670930951e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.20486160000956 lags = 1.56042886364135e-08 wags = -5.47752174539625e-08 pags = 8.72921955461756e-14   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.01403882011972+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.29606192622867e-07 wnfactor = -5.23018301329058e-08 pnfactor = 9.81789585875335e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -2.37230925107352 lpclm = 3.31327577293647e-06 wpclm = 3.03615475662011e-06 ppclm = -2.95861610764981e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -3.4566298065355e-06 lalpha0 = 2.57149637388823e-11 walpha0 = 5.58854999571259e-12 palpha0 = -2.38947528466507e-18   alpha1 = 0.0   beta0 = 20.4801076952924 lbeta0 = 1.32262083239532e-05 wbeta0 = 3.45922731795792e-06 pbeta0 = -3.04977933569516e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16473.456 lat = 0.006635672145984   ute = -0.863282674546883 lute = -7.10978310399278e-07 wute = -3.340527034145e-07 pute = 7.50270477982919e-13   ua1 = 3.0044e-9   ub1 = -3.04349011428923e-18 lub1 = -1.33409852530928e-24 wub1 = -9.87620992379907e-25 pub1 = 1.85834321361776e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.61 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.732619054637311+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.89845342572435e-08 wvth0 = 5.376755191693e-08 pvth0 = -3.66498990184482e-14   k1 = 0.88325   k2 = -0.0417049113707272 lk2 = 1.51815410698971e-08 wk2 = 5.53357264884414e-09 pk2 = -3.77188232606751e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4542.95159768406 lvsat = 0.0799288748435611 wvsat = 0.0487998380645189 pvsat = -3.32637264189465e-8   ua = -1.70291217752384e-10 lua = 2.03392123774639e-17 wua = -5.76605727063456e-18 pua = 3.93035221372632e-24   ub = 2.13241513919421e-18 lub = -1.17428936779787e-25 wub = -6.71814759440126e-25 pub = 4.57933125365728e-31   uc = 2.2391553446979e-10 luc = -1.0777246900185e-16 wuc = -2.17800805348183e-16 puc = 1.48460869754314e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0478549816675945 lu0 = -4.85780278517246e-09 wu0 = -3.21201630766237e-09 pu0 = 2.1894259478898e-15   a0 = 1.07852668459921 la0 = 2.97693040165296e-08 wa0 = -1.29357952766084e-07 pa0 = 8.81750374916621e-14   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.434927406112208 lags = -1.87230008392701e-07 wags = 1.95001959654669e-07 pags = -1.3292035577117e-13   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.62124243596103+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.1669724032127e-07 wnfactor = 2.60338911382402e-07 pnfactor = -1.77456374199055e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.60588526628508 lpclm = -1.0756797285695e-06 wpclm = -1.4091638632114e-06 ppclm = 9.60536819063963e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8646257938378e-06 lalpha0 = 2.01419172363916e-11 walpha0 = 1.2687957896775e-11 palpha0 = -8.64856886892612e-18   alpha1 = 0.0   beta0 = 30.44470996 lbeta0 = 4.44105624170546e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37954636 lkt1 = 6.00954836496017e-9   kt2 = -0.019151   at = 6959.10000000003 lat = 0.0150238709124   ute = -3.11005569428047 lute = 1.26985766762656e-06 wute = 2.27878794377687e-06 pute = -1.55330389884429e-12   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -1.39479310625539e-17 lub1 = 8.27964917455497e-24 wub1 = 4.93810496189954e-24 pub1 = -3.36599011380935e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.62 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.757917533840001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.17401800874378e-8   k1 = 0.88325   k2 = -0.0178715250696 lk2 = -1.06415303485813e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 128027.000392 lvsat = -0.00424229824040123   ua = -1.44942210792e-10 lua = 3.06041666901581e-18   ub = 1.711994052e-19 lub = 1.21940631127709e-24   uc = 8.143127184e-11 luc = -1.06500661599303e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.031222731904 lu0 = 6.47933741468506e-9   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.1791973824+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.63624937549606e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.704885509999999 lpclm = 1.18106082029436e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 6.309180502e-05 lalpha0 = -2.09110963026127e-11   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000007 lat = 0.015430120515312   ute = -1.12187464 lute = -8.535811348896e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.63 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.748192179871355+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.64242606714797e-08 wvth0 = 4.17070611337957e-08 pvth0 = -2.00876220962366e-14   k1 = 0.88325   k2 = 0.0349270468049523 lk2 = -2.649384599823e-08 wk2 = -2.63642172421759e-08 pk2 = 1.26979561356526e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 113908.410378837 lvsat = 0.00255772297917867 wvsat = -0.0265907436429618 pvsat = 1.28070594052215e-8   ua = -5.58004205498155e-11 lua = -3.98734786160691e-17 wua = -7.95624139357012e-17 pua = 3.83201227983354e-23   ub = 1.60399952048707e-18 lub = 5.29318194950688e-25 wub = 8.47432796904729e-25 pub = -4.08154142570007e-31   uc = -1.02323224239579e-10 luc = 7.78527143138541e-17 wuc = 1.88559968399337e-16 puc = -9.08172689399832e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0328342225358783 lu0 = 5.70318551270972e-09 wu0 = 7.03931265141173e-09 pu0 = -3.39038638817535e-15   a0 = 1.1222   keta = -0.01066   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.689623884229404+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.21712838152879e-08 wnfactor = 9.42752372088715e-08 pnfactor = -4.5406348148333e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.5123665 lpclm = -8.50119568794001e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.955060288e-05 lalpha0 = -9.57280586871168e-12   alpha1 = 0.0   beta0 = 36.96   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.447057199999999 lkt1 = 3.67619272992001e-8   kt2 = -0.019151   at = -63667.070749655 lat = 0.0491591756875809 wat = 0.0826356157770419 pat = -3.98002874403914e-8   ute = -0.239122371498592 lute = -5.10523385080904e-07 wute = -1.4791623320385e-06 pute = 7.12417828953696e-13   ua1 = -1.776800572e-09 lua1 = 1.82467826149579e-15   ub1 = 1.92300317206582e-17 lub1 = -1.0129398321011e-23 wub1 = -1.89224547110779e-23 pub1 = 9.11373539722473e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.64 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.7328083932272+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.50962870646259e-8   k1 = 0.88325   k2 = -0.04434110208 wk2 = 7.90009057915263e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 139932.9688 wvsat = -0.0250322637537104   ua = -1.634473084208e-10 wua = 1.46046034968208e-17   ub = 1.5945968728e-19 wub = 1.47371137370582e-24   uc = 4.1443099808e-11 wuc = 1.00037193496479e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0346737890268 wu0 = 3.16084001994673e-9   a0 = 1.9166505784264 wa0 = -7.12828617763881e-7   keta = -0.025911781888 wketa = 3.6377161271447e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.219567414024 wags = -3.81386058860429e-8   b0 = 5.6910853536e-07 wb0 = -4.78782233703995e-13   b1 = -1.87957198056e-09 wb1 = 1.6783788366169e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.05427077328+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.87985860065618e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.14243742536 wpclm = -1.88828240607461e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.7884966168e-05 walpha0 = -6.31318284944496e-12   alpha1 = 0.0   beta0 = 22.43957568 wbeta0 = 4.04190680793854e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.397873664 wkt1 = 4.59307591811182e-9   kt2 = -0.019151   at = 381464.88 wat = -0.20668841631504   ute = -1.261285952 wute = 8.26753665260158e-8   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.65 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.684927712800005+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.5194625968582e-07 wvth0 = 1.07851723697533e-07 pvth0 = -8.50048028156531e-13   k1 = 0.88325   k2 = -0.0501519052674503 lk2 = 1.15528273840525e-07 wk2 = 1.30888937718118e-08 pk2 = -1.03161896352088e-13   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 158345.106806746 lvsat = -0.366063425831897 wvsat = -0.0414735296839386 pvsat = 3.26879264603999e-7   ua = -1.74189524057507e-10 lua = 2.13572821122511e-16 wua = 2.4196950887343e-17 pua = -1.90711559203915e-22   ub = -9.24508485225435e-19 lub = 2.15510606413383e-23 wub = 2.44164942508993e-24 pub = -1.92441920081681e-29   uc = 3.40850013531938e-11 luc = 1.46291035130619e-16 wuc = 1.65741922296548e-17 puc = -1.30631750148167e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0323488765363793 lu0 = 4.62230638663974e-08 wu0 = 5.23688922756779e-09 pu0 = -4.12752546640105e-14   a0 = 2.44096188381049 la0 = -1.04241665243314e-05 wa0 = -1.18101659239705e-06 pa0 = 9.30834289123393e-12   keta = -0.0285874540533841 lketa = 5.31967400474976e-08 wketa = 6.02697899260173e-09 pketa = -4.75024545993335e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.247619742086205 lags = -5.57726175485349e-07 wags = -6.31881566478137e-08 pags = 4.98026050209047e-13   b0 = 9.21270235511054e-07 lb0 = -7.0015507355444e-12 wb0 = -7.9324784114748e-13 pb0 = 6.25209074171026e-18   b1 = -3.11408049610775e-09 lb1 = 2.45440489450207e-14 wb1 = 2.78074309164338e-15 pb1 = -2.19168048578478e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.07545317792262+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.21140858709355e-07 wnfactor = -4.77135836914307e-08 pnfactor = 3.76061098911392e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 4.53133763024872 lpclm = -2.7613608313923e-05 wpclm = -3.12851195523164e-06 ppclm = 2.46577924527841e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.25285411570409e-05 lalpha0 = -9.23218676708153e-11 walpha0 = -1.04597002845089e-11 palpha0 = 8.24395503115959e-17   alpha1 = 0.0   beta0 = 19.4666066073511 lbeta0 = 5.91074889416641e-05 wbeta0 = 6.69664332511302e-06 pbeta0 = -5.27805051103705e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.401252037946192 lkt1 = 6.71676010700713e-08 wkt1 = 7.60982196035567e-09 pkt1 = -5.99778467163299e-14   kt2 = -0.019151   at = 533491.70757864 lat = -3.02254204815328 wat = -0.342441988216007 pat = 2.69900310223486e-6   ute = -1.32209668303146 lute = 1.20901681926131e-06 wute = 1.36976795286403e-07 pute = -1.07960124089394e-12   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.66 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.851833923006003+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.63547735297337e-07 wvth0 = -4.73426398312897e-08 pvth0 = 3.73137454429327e-13   k1 = 0.88325   k2 = -0.0340985024036284 lk2 = -1.09988040934759e-08 wk2 = -3.0435732141556e-09 pk2 = 2.39883362133243e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 84696.5547797609 lvsat = 0.214407653171865 wvsat = 0.0242915340369744 pvsat = -1.91457029161043e-7   ua = -1.450651095879e-10 lua = -1.59752124400619e-17 wua = -5.27104002791305e-18 pua = 4.15444188414405e-23   ub = 1.5381246276963e-18 lub = 2.14148284374229e-24 wub = -2.25688408433431e-25 pub = 1.77879388469163e-30   uc = 6.35173951724186e-11 luc = -8.56843795611601e-17 wuc = -9.70769929037251e-18 puc = 7.65125522041744e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0364725427431893 lu0 = 1.37218278388208e-08 wu0 = 2.60632560148996e-10 pu0 = -2.05421096884253e-15   a0 = 0.377028673975018 la0 = 5.84300376390344e-06 wa0 = 6.70317081716441e-07 pa0 = -5.28319524267125e-12   keta = -0.0178847653918478 lketa = -3.11579562040581e-08 wketa = -3.53007246922636e-09 pketa = 2.78227462560634e-14   a1 = 0.0   a2 = 0.65972622   ags = -0.0529464369725641 lags = 1.81122704176669e-06 wags = 1.5811560076966e-07 pags = -1.24620961118778e-12   b0 = -4.87376565093162e-07 lb0 = 4.10089059938261e-12 wb0 = 4.6461458862646e-13 pb0 = -3.6619230678435e-18   b1 = 1.82395356608325e-09 lb1 = -1.43757380887701e-14 wb1 = -1.62871392846256e-15 pb1 = 1.2836930332272e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.06472560392893+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.36590025327975e-07 wnfactor = -1.96337995289679e-08 pnfactor = 1.54746461184292e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.02426318930617 lpclm = 1.61736151071103e-05 wpclm = 1.83240624139646e-06 ppclm = -1.4442358998815e-11   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 5.55446221972681e-05 lalpha0 = -1.94909880576388e-10 walpha0 = -1.41849187289304e-11 palpha0 = 1.11800366111012e-16   alpha1 = 0.0   beta0 = 27.4625438766672 lbeta0 = -3.91357809391944e-06 wbeta0 = -1.41737758234089e-06 pbeta0 = 1.11712541785709e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.394670818 lkt1 = 1.52968210182501e-8   kt2 = -0.019151   at = 306659.56838576 lat = -1.23473369393367 wat = -0.0445716220861914 pat = 3.51297301212922e-7   ute = -1.07885375890563 lute = -7.08135368274052e-07 wute = -8.02289197551443e-08 pute = 6.3233514218326e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.67 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.752538367036567+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.18814693936418e-08 wvth0 = 5.28253454515432e-08 pvth0 = -1.56782032919874e-14   k1 = 0.88325   k2 = -0.0427866410751313 lk2 = 2.27253877468219e-08 wk2 = 4.97636950161079e-09 pk2 = -7.14216215013198e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 170514.070479054 lvsat = -0.118704705197078 wvsat = -0.0507436923235118 pvsat = 9.98024067479698e-8   ua = -1.44731305655129e-10 lua = -1.72709178024483e-17 wua = 3.24565196505143e-18 pua = 8.48572060063813e-24   ub = 2.34395666459811e-18 lub = -9.86463800649128e-25 wub = 4.10562624792613e-25 pub = -6.9090103091578e-31   uc = -2.78370155149874e-12 luc = 1.71672344321879e-16 wuc = 3.84396950981485e-17 puc = -1.10378107160507e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.038548734424831 lu0 = 5.66280746445969e-09 wu0 = 7.64068639524647e-10 pu0 = -4.0083665782458e-15   a0 = 1.54767815256893 la0 = 1.29896860441207e-06 wa0 = -3.94138140923755e-07 pa0 = -1.15136753008305e-12   keta = -0.025911781888 wketa = 3.6377161271447e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.505854964391655 lags = -3.5783659461911e-07 wags = -2.2220947669533e-07 pags = 2.30073901203114e-13   b0 = 8.31962168707864e-07 lb0 = -1.02030212593387e-12 wb0 = -7.13499488431037e-13 pb0 = 9.1108694576966e-19   b1 = -2.20336631027824e-09 lb1 = 1.25685172683019e-15 wb1 = 1.96751357369344e-15 pb1 = -1.12231580428683e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.2147199744211+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.18813573627748e-07 wnfactor = -1.44385462154932e-07 pnfactor = 6.38987005893092e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.14243742536 wpclm = -1.88828240607461e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.76950430657233e-05 lalpha0 = -8.68079516345343e-11 walpha0 = 2.38509728548672e-13 palpha0 = 5.58138669670369e-17   alpha1 = 0.0   beta0 = 27.5318041993475 lbeta0 = -4.18242145580719e-06 wbeta0 = -7.43238592594808e-07 pbeta0 = 8.55449200696881e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284644e-8   kt2 = -0.019151   at = -41012.7967715199 lat = 0.114803874865976 wat = 0.0891432441723829 pat = -1.67735137391546e-7   ute = -1.34839248218874 lute = 3.38115843415685e-07 wute = 1.60457839510289e-07 pute = -3.01923247304784e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.68 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.723452785525398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.66099466459894e-08 wvth0 = 6.36296780882257e-08 pvth0 = -3.60080245371428e-14   k1 = 0.88325   k2 = -0.032704215138543 lk2 = 3.75393213720373e-09 wk2 = -2.00361210161787e-09 pk2 = 5.99162251384066e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 104782.513077981 lvsat = 0.00497815954484848 wvsat = 0.00654843009320361 pvsat = -8.000513307729e-9   ua = -1.38337225036031e-10 lua = -2.93022500822448e-17 wua = -3.42544785664408e-18 pua = 2.10383021847339e-23   ub = 1.91785045561191e-18 lub = -1.84687017997176e-25 wub = -1.29863393889896e-26 pub = 1.06063947851034e-31   uc = 1.49745200460087e-10 luc = -1.15331528743592e-16 wuc = -5.96299826814163e-17 puc = 7.41533290579224e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0399340311695974 lu0 = 3.05618323882433e-09 wu0 = -1.09728565963604e-09 pu0 = -5.05975320190249e-16   a0 = 3.35644872481106 la0 = -2.10447922005931e-06 wa0 = -1.97958891481707e-06 pa0 = 1.83187372230247e-12   keta = -0.0393583018646088 lketa = 2.53014560627062e-08 wketa = 6.84485762261604e-09 pketa = -6.03467289497272e-15   a1 = 0.0   a2 = 0.65972622   ags = 0.100494270669495 lags = 4.0490467967348e-07 wags = 3.84204242188826e-08 pags = -2.60336703033501e-13   b0 = 1.00701994101352e-08 lb0 = 5.26199391607629e-13 wb0 = 2.04155206891245e-14 pb0 = -4.69873956331165e-19   b1 = -1.13217150693529e-09 lb1 = -7.58746978152827e-16 wb1 = 1.01098160448992e-15 pb1 = 6.77529184117392e-22   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.669904763533701+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.0633034052558e-07 wnfactor = 2.54995428768036e-07 pnfactor = -1.12502456179637e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 5.58950476353275 lpclm = -4.60448999793002e-06 wpclm = -4.07341076223468e-06 ppclm = 4.1116161795716e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -6.21733378842869e-05 lalpha0 = 8.22916292227191e-11 walpha0 = 5.80201042074054e-11 palpha0 = -5.29100613417811e-17   alpha1 = 0.0   beta0 = 16.3402039186363 lbeta0 = 1.68760965299891e-05 wbeta0 = 7.15598751455313e-06 pbeta0 = -6.30897620838058e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16473.456 lat = 0.006635672145984   ute = -1.70854925331219 lute = 1.01579978960533e-06 wute = 4.20734850226607e-07 pute = -7.91669840640993e-13   ua1 = 3.0044e-9   ub1 = -4.49029386827594e-18 lub1 = 1.38825950312728e-24 wub1 = 3.04313994172565e-25 pub1 = -5.72608166738888e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.69 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.730143796011188+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.07109109253403e-08 wvth0 = 5.59778539091942e-08 pvth0 = -2.92619008752404e-14   k1 = 0.88325   k2 = -0.0455205002080528 lk2 = 1.5053230440746e-08 wk2 = 8.94073322584467e-09 pk2 = -3.65730632328212e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 104013.373880261 lvsat = 0.0056562603505701 wvsat = -0.0400230712760856 pvsat = 3.30585988734859e-8   ua = -2.58221007287543e-10 lua = 7.63916081668489e-17 wua = 7.27515517331021e-17 pua = -4.61220830255716e-23   ub = 1.16653579743166e-18 lub = 4.77699031982232e-25 wub = 1.90674925821481e-25 pub = -7.34911553640629e-32   uc = -1.91367707927722e-10 luc = 1.85405891355802e-16 wuc = 1.53029688216615e-16 puc = -1.13335092553934e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0498099872277807 lu0 = -5.65081515648811e-09 wu0 = -4.95775416267502e-09 pu0 = 2.89755268895497e-15   a0 = 0.448774443441046 la0 = 4.59031102670622e-07 wa0 = 4.32984348994034e-07 pa0 = -2.95137719710899e-13   keta = 0.0435338890098769 lketa = -4.77792835311119e-08 wketa = -4.83928667424817e-08 pketa = 4.26648934633746e-14   a1 = 0.0   a2 = 0.65972622   ags = 1.92135938744726 lags = -1.200435558422e-06 wags = -1.13231936953431e-06 pags = 7.71829645771891e-13   b0 = 2.56314661773392e-06 lb0 = -1.72468468953768e-12 wb0 = -2.25937449166444e-12 pb0 = 1.54007099100018e-18   b1 = -8.78455068420613e-09 lb1 = 5.98786599017953e-15 wb1 = 7.84423480986734e-15 pb1 = -5.34691283885874e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.171549521076452+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.4569826306462e-07 wnfactor = 6.61895797271905e-07 pnfactor = -4.71240469465913e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.21003224679822 lpclm = 1.39022661371013e-06 wpclm = 1.99829020743645e-06 ppclm = -1.24141397652538e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.58798335653201e-05 lalpha0 = 4.66078335857344e-12 walpha0 = -7.86365600443224e-12 palpha0 = 5.17543347634258e-18   alpha1 = 0.0   beta0 = 30.4447099600001 lbeta0 = 4.44105624170541e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.379546360000001 lkt1 = 6.00954836496102e-9   kt2 = -0.019151   at = 6959.10000000003 lat = 0.0150238709123999   ute = 1.79774757856093 lute = -2.07547772405996e-06 wute = -2.10367425113304e-06 pute = 1.43394010184532e-12   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -6.71391229262028e-18 lub1 = 3.34868155629251e-24 wub1 = -1.52156997086283e-24 pub1 = 1.03715686865905e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.70 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.707289563462806+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.6289178582689e-08 wvth0 = 4.52086511720791e-08 pvth0 = -2.19212245983233e-14   k1 = 0.88325   k2 = -0.0045704019786357 lk2 = -1.28598307159609e-08 wk2 = -1.18773442730613e-08 pk2 = 1.05330447507622e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 156111.325791444 lvsat = -0.029855579198362 wvsat = -0.0250781230400372 pvsat = 2.28715841376587e-8   ua = -1.66243585996284e-10 lua = 1.36964866275603e-17 wua = 1.90212333996669e-17 pua = -9.497563758042e-24   ub = -2.61678913501118e-18 lub = 3.05654950563284e-24 wub = 2.48955667088989e-24 pub = -1.64049171254552e-30   uc = 1.66187950969616e-10 luc = -5.8316917752344e-17 wuc = -7.56841546822238e-17 puc = 4.25644964642586e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0261138568542866 lu0 = 1.05013203667789e-08 wu0 = 4.56201084664212e-09 pu0 = -3.59146185293587e-15   a0 = 1.1222   keta = -0.0265611228896 wketa = 1.41990348932514e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.49359792712893+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.55457524243369e-07 wnfactor = -2.8074648162006e-07 pnfactor = 1.71298442948889e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -5.35934979775432 lpclm = 4.21855083187364e-06 wpclm = 4.15624112146452e-06 ppclm = -2.71235100575981e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 6.2286656440949e-05 lalpha0 = -2.01554177590788e-11 walpha0 = 7.18963864852254e-13 palpha0 = -6.7478920087702e-19   alpha1 = 0.0   beta0 = 34.7303636211264 lbeta0 = 1.51980042274987e-06 wbeta0 = 1.9909716416062e-06 pbeta0 = -1.3571179458979e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000001 lat = 0.015430120515312   ute = -1.12187464 lute = -8.53581134889591e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.71 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.744104524436381+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.85577680392208e-08 wvth0 = 4.53571657556999e-08 pvth0 = -2.19927545683194e-14   k1 = 0.88325   k2 = -0.00418820803014391 lk2 = -1.30439090805367e-08 wk2 = 8.564062484862e-09 pk2 = 6.87727365503006e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 34124.1556362824 lvsat = 0.0288978334864898 wvsat = 0.0446532449034402 pvsat = -1.0713552993166e-8   ua = -6.88370904744419e-11 lua = -3.32179882495977e-17 wua = -6.7921215233147e-17 pua = 3.23770494316717e-23   ub = 9.80793366971888e-18 lub = -2.92764428714613e-24 wub = -6.47833583312501e-24 pub = 2.67876816151821e-30   uc = -4.14867862194393e-11 luc = 4.17067119684439e-17 wuc = 1.34235584377749e-16 puc = -5.85404069776304e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.041302324158317 lu0 = 3.18600772833482e-09 wu0 = -5.22346437158145e-10 pu0 = -1.14265234819549e-15   a0 = 1.1222   keta = -0.0872455322405538 lketa = 2.9227796182156e-08 wketa = 6.83876636984604e-08 pketa = -2.60991944232257e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.1755583034529+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.02278192054537e-07 wnfactor = -3.39643789912098e-07 pnfactor = 1.99665506925434e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 11.4696909988244 lpclm = -3.88692106122737e-06 wpclm = -7.10555656982128e-06 ppclm = 2.71173618708031e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.32295029051414e-05 lalpha0 = -1.09768065587065e-11 walpha0 = -3.28510320865025e-12 palpha0 = 1.25371364813644e-18   alpha1 = 0.0   beta0 = 41.4192727577471 lbeta0 = -1.7018190181756e-06 wbeta0 = -3.98194328321241e-06 pbeta0 = 1.51965290683205e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4470572 lkt1 = 3.67619272992003e-8   kt2 = -0.019151   at = 28874.36544 lat = 0.0045878885269402   ute = -1.895597068 lute = 2.87294461843246e-7   ua1 = -1.77680057200001e-09 lua1 = 1.82467826149579e-15   ub1 = -4.31535116948764e-18 lub1 = 1.21090571266735e-24 wub1 = 2.10258330374096e-24 pub1 = -1.01267981208058e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.72 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.8340534+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}   k1 = 0.88325   k2 = -0.032054   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 101000.0   ua = -1.407326e-10   ub = 2.45154e-18   uc = 5.7002e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03958988   a0 = 0.80798   keta = -0.020254   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -1.75547e-7   b1 = 7.3083e-10   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00948+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.20557   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8066e-5   alpha1 = 0.0   beta0 = 28.726   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.39073   kt2 = -0.019151   at = 60000.0   ute = -1.1327   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.73 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.852670743756203+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.70143251847638e-7   k1 = 0.88325   k2 = -0.02979459768 lk2 = -4.49206145037955e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 93840.8473 lvsat = 0.142335668049817   ua = -1.365557270018e-10 lua = -8.30430685684455e-17   ub = 2.87301705313e-18 lub = -8.37965335268329e-24   uc = 5.98630338679998e-11 luc = -5.68820339472484e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0404938708090501 lu0 = -1.79728162128782e-8   a0 = 0.604113143461902 la0 = 4.05320663415473e-6   keta = -0.019213624048 lketa = -2.06843759808174e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.149342472579 lags = 2.1685948984434e-7   b0 = -3.1247728944e-07 lb0 = 2.72239817202073e-12   b1 = 1.21084133649e-09 lb1 = -9.5434106679677e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.00124369038+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.63751309848148e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.33447313069 lpclm = 1.0736940948679e-05 ppclm = -3.23117426778526e-27   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.6260448553e-05 lalpha0 = 3.58973166485275e-11   alpha1 = 0.0   beta0 = 29.8819732799999 lbeta0 = -2.29826399786867e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.389416393999999 lkt1 = -2.61166363394242e-8   kt2 = -0.019151   at = 887.730000000214 lat = 1.17524863527372   ute = -1.109055092 lute = -4.70099454109499e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.74 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.778201368731402+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.16797255245328e-7   k1 = 0.88325   k2 = -0.0388322069599999 lk2 = 2.63105321513865e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 122477.4581 lvsat = -0.0833676745494536   ua = -1.532632189946e-10 lua = 4.86393017917233e-17   ub = 1.18710884061001e-18 lub = 4.90806150780993e-24   uc = 4.84188983960002e-11 luc = 3.33164761777442e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.03687790757285 lu0 = 1.0526889804233e-8   a0 = 1.41958056961429 la0 = -2.37401078863538e-6   keta = -0.023375127856 lketa = 1.21150822464524e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.192972582263001 lags = -1.27017153325026e-7   b0 = 2.3524386832e-07 lb0 = -1.59454062294217e-12 wb0 = 1.0097419586829e-28 pb0 = 3.85185988877447e-34   b1 = -7.09204009470001e-10 lb1 = 5.58968785238309e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.03418892886+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.59110677844116e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.82569939207 lpclm = -6.28875257291703e-6   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.3482654341e-05 lalpha0 = -2.10254804895817e-11   alpha1 = 0.0   beta0 = 25.25808016 lbeta0 = 1.34612024960583e-5   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.394670818 lkt1 = 1.52968210182433e-8   kt2 = -0.019151   at = 237336.81 lat = -0.688356945821161   ute = -1.203634724 lute = 2.7534277832846e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.75 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.8346982366572+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.50302118270864e-9   k1 = 0.88325   k2 = -0.0350468361398 lk2 = 1.16171005023488e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 91591.8200000003 lvsat = 0.0365191301824801   ua = -1.396833056846e-10 lua = -4.07297858925198e-18   ub = 2.98250945466001e-18 lub = -2.06103015010864e-24   uc = 5.7002e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0397370992006401 lu0 = -5.7145134909524e-10   a0 = 0.93467055188 la0 = -4.91766607037276e-7   keta = -0.020254   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -2.77751822612e-07 lb0 = 3.96721918824354e-13   b1 = 8.56730264759999e-10 lb1 = -4.88699000101946e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.990155598280001+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.5010293394814e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.20557   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8066e-5   alpha1 = 0.0   beta0 = 26.3758366359999 lbeta0 = 9.12247871958337e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284644e-8   kt2 = -0.019151   at = 97632.7200000002 lat = -0.14607652072992   ute = -1.098830552 lute = -1.31468868656922e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.76 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.822416758426002+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.06062503903364e-8   k1 = 0.88325   k2 = -0.0358204561708 lk2 = 1.30727718029993e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 114967.362 lvsat = -0.0074651311642322   ua = -1.436648636324e-10 lua = 3.41886418141459e-18   ub = 1.89765265204e-18 lub = -1.9724535453938e-26   uc = 5.7002e-11   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0382274101156 lu0 = 2.2692339821229e-9   a0 = 0.277571232320003 la0 = 7.44655128222325e-7   keta = -0.028712415784 lketa = 1.59156596421426e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 4.18226944240003e-08 lb0 = -2.04600997113197e-13 pb0 = -9.62964972193618e-35   b1 = 4.40219853759998e-10 lb1 = 2.95021983610449e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.06650209768+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.86460283502034e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.74591802028 lpclm = 1.79035411252758e-06 wpclm = 4.2351647362715e-22 ppclm = 4.03896783473158e-28   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 2.8066e-5   alpha1 = 0.0   beta0 = 27.4699939119999 lbeta0 = 7.06367299939988e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16473.4560000001 lat = 0.00663567214598404   ute = -1.0541754836 lute = -2.15493452940832e-7   ua1 = 3.0044e-9   ub1 = -4.0169908e-18 lub1 = 4.97675410948811e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.77 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.81720679843+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.51995386813753e-8   k1 = 0.88325   k2 = -0.0316148746060001 lk2 = 9.36497969453545e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 41765.0290799998 lvsat = 0.0570726808220261   ua = -1.45069679e-10 lua = 4.65739998284389e-18   ub = 1.46309471080001e-18 lub = 3.63397389629133e-25   uc = 4.66411328000002e-11 luc = 9.13451351473958e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0420991349439999 lu0 = -1.1442180086882e-9   a0 = 1.1222   keta = -0.031732095304 lketa = 1.85779178154373e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -9.50884612399999e-07 lb0 = 6.70605502045887e-13   b1 = 3.415678273e-09 lb1 = -2.32824927529463e-15   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.2010036958+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.87227479310328e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.897931582 lpclm = -5.40558875428153e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.36493985999999e-05 lalpha0 = 1.27101947918904e-11   alpha1 = 0.0   beta0 = 30.4447099600002 lbeta0 = 4.44105624170551e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.379546359999999 lkt1 = 6.00954836495848e-9   kt2 = -0.019151   at = 6959.10000000009 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397724e-7   ua1 = 6.387700286e-09 lua1 = -2.98283933094789e-15   ub1 = -9.08042763399999e-18 lub1 = 4.96178360752923e-24   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.78 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.777603100540006+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.21948448963197e-8   k1 = 0.88325   k2 = -0.023043372644 lk2 = 3.52233538316559e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 117107.031514001 lvsat = 0.00571685965092295   ua = -1.36659642100001e-10 lua = -1.07518392952452e-18   ub = 1.25524709580001e-18 lub = 5.05073806527271e-25   uc = 4.84755114600001e-11 luc = 7.88413498245148e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0332092049900001 lu0 = 4.91547828543631e-9   a0 = 1.1222   keta = -0.0044772   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.0569496832+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.90350783777114e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 1.1049   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 6.34048692399998e-05 lalpha0 = -2.12049251932767e-11   alpha1 = 0.0   beta0 = 37.8269448000003 lbeta0 = -5.90940785692804e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000024 lat = 0.015430120515312   ute = -1.12187464 lute = -8.53581134889566e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.79 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.814649047959996+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.43521829647371e-8   k1 = 0.88325   k2 = 0.00913157721999991 lk2 = -1.19742787695319e-8   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 103573.862931999 lvsat = 0.0122349208340831   ua = -1.74475740639999e-10 lua = 1.71384105068869e-17   ub = -2.67896840400005e-19 lub = 1.2386747593829e-24   uc = 1.6729136784e-10 luc = -4.93418588209864e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0404899127143996 lu0 = 1.40882733988747e-9   a0 = 1.1222   keta = 0.019118590608 lketa = -1.13645822052747e-8   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.647306396000005+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.08263875896139e-7   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 0.418336835999995 lpclm = 3.30673536056306e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 3.81201439599999e-05 lalpha0 = -9.0268912483186e-12   alpha1 = 0.0   beta0 = 35.2261103999999 lbeta0 = 6.61714691385607e-7   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.4470572 lkt1 = 3.67619272991999e-8   kt2 = -0.019151   at = 28874.3654400003 lat = 0.00458788852694014   ute = -1.895597068 lute = 2.87294461843251e-7   ua1 = -1.77680057199999e-09 lua1 = 1.8246782614958e-15   ub1 = -1.045179084e-18 lub1 = -3.64126889898572e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.80 nmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.837534387125714+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.06407916408921e-9   k1 = 0.88325   k2 = -0.0352618195 wk2 = 1.902102235081e-9   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 70039.5121428571 wvsat = 0.0183582689587957   ua = -3.0922762241e-10 wua = 9.99104714981888e-17   ub = 2.92570043038571e-18 wub = -2.81157220480653e-25   uc = 3.33993782642857e-11 wuc = 1.39953633791657e-17   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0381029718337143 wu0 = 8.81674092464449e-10   a0 = 0.477116331571429 wa0 = 1.96188259104069e-7   keta = -0.0262493811142857 wketa = 3.55500919476463e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -3.59939618185714e-07 wb0 = 1.09337078094165e-13   b1 = 1.24144333114286e-09 wb1 = -3.02772259607806e-16   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.871443167857143+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor = 8.18500439137643e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.123482982857143 wpclm = 1.95114598609006e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.76087319714286e-05 walpha0 = 6.20072073568566e-12   alpha1 = 0.0   beta0 = 33.7087384428571 wbeta0 = -2.95455462159969e-6   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.394083121428571 wkt1 = 1.98826017604285e-9   kt2 = -0.019151   at = -163541.428571429 wat = 0.132550678402857   ute = -1.23754093 wute = 6.216626817094e-8   ua1 = 3.0044e-9   ub1 = -4.08803568428571e-18 wub1 = 1.98958568282688e-25   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.81 nmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.881021804567237+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.64601004152421e-07 wvth0 = -1.68109883163913e-08 pvth0 = 2.93192679891139e-13   k1 = 0.88325   k2 = -0.0295607467167887 lk2 = -1.13346653885314e-07 wk2 = -1.38663799443858e-10 pk2 = 4.05737674595866e-14   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 54878.5233332621 lvsat = 0.301425260912441 wvsat = 0.0231030216946689 pvsat = -9.43334468046359e-8   ua = -2.97645453854742e-10 lua = -2.30272459306279e-16 wua = 9.5519442255267e-17 pua = 8.7300845073127e-23   ub = 4.12936503847608e-18 lub = -2.39308216041352e-23 wub = -7.44961588694838e-25 pub = 9.22118962404442e-30   uc = 3.94582101225055e-11 luc = -1.2045948959033e-16 wuc = 1.20992034784809e-17 puc = 3.76987609432104e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0405088485514629 lu0 = -4.78327651631529e-08 wu0 = -8.88117218567351e-12 pu0 = 1.77056956096573e-14   a0 = -0.100746581020862 la0 = 1.14888600860597e-05 wa0 = 4.1795221250985e-07 pa0 = -4.40903019953469e-12   keta = -0.0240461695294785 lketa = -4.38034507601198e-08 wketa = 2.86549650360654e-09 pketa = 1.37086403429856e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.137151051269638 lags = 4.59244890639716e-07 wags = 7.22900079675658e-09 pags = -1.43724362484824e-13   b0 = -6.39089697489186e-07 lb0 = 5.54996026608276e-12 wb0 = 1.93667440252029e-13 pb0 = -1.67662556417083e-18   b1 = 1.98089768593487e-09 lb1 = -1.47015623205897e-14 wb1 = -4.56611072854133e-16 pb1 = 3.05856728763544e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.832102473286359+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.82157369443496e-07 wnfactor = 1.00293637805411e-07 pnfactor = -3.66688820285542e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.26713617817029 lpclm = 2.27376965394529e-05 wpclm = 5.53030015307818e-07 ppclm = -7.1159440335941e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 1.57532863084499e-06 lalpha0 = 3.18770289058666e-10 walpha0 = 1.46372393388012e-11 palpha0 = -1.67731791974371e-16   alpha1 = 0.0   beta0 = 36.8989399668652 lbeta0 = -6.34264254669733e-05 wbeta0 = -4.16076653271021e-06 pbeta0 = 2.39814661555638e-11   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.402312989687721 lkt1 = 1.63623245056373e-07 wkt1 = 7.64713958579988e-09 pkt1 = -1.12507780592685e-13   kt2 = -0.019151   at = -338643.616490329 lat = 3.48131796300717 wat = 0.201327828152212 pat = -1.36740225643417e-6   ute = -1.24465537365065 lute = 1.41446779004639e-07 wute = 8.04052718070035e-08 pute = -3.62621231294886e-13   ua1 = 3.0044e-9   ub1 = -4.30841652833162e-18 lub1 = 4.38153172269356e-24 wub1 = 3.29635152806463e-25 pub1 = -2.59806428722492e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.82 nmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.726199639004576+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.55650949544216e-07 wvth0 = 3.08348416553583e-08 pvth0 = -8.23344088640818e-14   k1 = 0.88325   k2 = -0.0491555001298508 lk2 = 4.10920600261988e-08 wk2 = 6.12127927140837e-09 pk2 = -8.76482520559299e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 109014.680146885 lvsat = -0.125256221531454 wvsat = 0.00798286188952316 pvsat = 2.48381490413542e-8   ua = -3.42400325490053e-10 lua = 1.22469148149961e-16 wua = 1.12150360393331e-16 pua = -4.37779980368882e-23   ub = -4.39617495552359e-19 lub = 1.20802356194345e-23 wub = 9.64580394838162e-25 pub = -4.25279801688069e-30   uc = -1.14731910817982e-11 luc = 2.80963275671954e-16 wuc = 3.55134935925763e-17 puc = -1.46844150934488e-22   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0321442752857377 lu0 = 1.80937566126245e-08 wu0 = 2.80684513370153e-09 pu0 = -4.48683420897036e-15   a0 = 1.99479801027627 la0 = -5.02745960431305e-06 wa0 = -3.41079783180042e-07 pa0 = 1.5733837028466e-12   keta = -0.039139041348598 lketa = 7.51530711128373e-08 wketa = 9.3473386167439e-09 pketa = -3.73788798022339e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.229546846191086 lags = -2.6898513286178e-07 wags = -2.16870023902697e-08 pags = 8.4181049210157e-14   b0 = 4.6147757367224e-07 lb0 = -3.1243103587249e-12 wb0 = -1.34147085458254e-13 pb0 = 9.07089202990257e-19   b1 = -2.39011316180685e-10 lb1 = 2.79495238720835e-15 wb1 = -2.78804519027446e-16 pb1 = 1.65716075195909e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.973889920672908+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.35359680226432e-07 wnfactor = 3.57547792966018e-08 pnfactor = 1.41982970336394e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 3.3074766030823 lpclm = -1.33177362433276e-05 wpclm = -8.78631651487429e-07 ppclm = 4.16789209923932e-12   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.09999160074472e-05 lalpha0 = 8.04004190609315e-12 walpha0 = -4.45742044321318e-12 palpha0 = -1.72346340286947e-17   alpha1 = 0.0   beta0 = 26.3768165289495 lbeta0 = 1.95051214177471e-05 wbeta0 = -6.63363679859526e-07 pbeta0 = -3.58379007596683e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.3726474158635 lkt1 = -7.01900095572666e-08 wkt1 = -1.30589524840547e-08 pkt1 = 5.0690100084396e-14   kt2 = -0.019151   at = 166531.182442557 lat = -0.500285918555027 wat = 0.0419847633052062 pat = -1.11518220185672e-7   ute = -1.31793618108844 lute = 7.19019429015391e-07 wute = 6.77759633922444e-08 pute = -2.63081619438018e-13   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.83 nmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.811405557147768+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.49125902665466e-08 wvth0 = 1.38115806565537e-08 pvth0 = -1.62563061337265e-14   k1 = 0.88325   k2 = -0.0379867622505514 lk2 = -2.26091500065312e-09 wk2 = 1.74325270677895e-09 pk2 = 8.22908031662897e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 54718.8670152571 lvsat = 0.0855003613695454 wvsat = 0.0218641124559271 pvsat = -2.90438128822199e-8   ua = -3.81686481962269e-10 lua = 2.74963707414148e-16 wua = 1.43497719399254e-16 pua = -1.65457035259204e-22   ub = 3.56793079754509e-18 lub = -3.47560810679107e-24 wub = -3.47130268634456e-25 pub = 8.3878531603851e-31   uc = 6.85816786261522e-11 luc = -2.97805885617357e-17 wuc = -6.86626307880598e-18 puc = 1.76586382323897e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0361169630743707 lu0 = 2.67322867550636e-09 wu0 = 2.1465886771604e-09 pu0 = -1.92395897802784e-15   a0 = 0.865941441560639 la0 = -6.45649308349974e-07 wa0 = 4.07534757967478e-08 pa0 = 9.12459788049744e-14   keta = -0.0197778567571429 wketa = -2.82332944998087e-10   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -5.8528109599214e-07 lb0 = 9.38825776756465e-13 wb0 = 1.82351942884941e-13 pb0 = -3.21444819391709e-19   b1 = 3.05937979223763e-09 lb1 = -1.00082012813081e-14 wb1 = -1.30607865851408e-15 pb1 = 5.64466503365944e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.80901884703009+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.04609814584181e-07 wnfactor = 1.07406485747645e-07 pnfactor = -1.36142872885406e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.123482982857143 wpclm = 1.95114598609006e-7   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.44098529982386e-05 lalpha0 = -5.19609227509454e-12 walpha0 = -9.69121838612957e-12 palpha0 = 3.08106448325549e-18   alpha1 = 0.0   beta0 = 30.2009815216103 lbeta0 = 4.66110491229501e-06 wbeta0 = -2.26815026108173e-06 pbeta0 = 2.64540729002218e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.407664724 lkt1 = 6.57344343284644e-8   kt2 = -0.019151   at = 54247.3971682857 lat = -0.0644411354181446 wat = 0.0257256742556477 pat = -4.84063548036998e-8   ute = -1.098830552 lute = -1.31468868656927e-7   ua1 = 3.0044e-9   ub1 = -3.7525e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.84 nmos  lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.826046789650981+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.6368798958693e-09 wvth0 = -2.15245605510253e-09 pvth0 = 1.37822000482471e-14   k1 = 0.88325   k2 = -0.0467435900369747 lk2 = 1.42162474080812e-08 wk2 = 6.4769596110192e-09 pk2 = -6.78033007838056e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 111565.454666516 lvsat = -0.0214642244322182 wvsat = 0.00201718816864818 pvsat = 8.30087434599859e-9   ua = -2.382423525515e-10 lua = 5.05406952618777e-18 wua = 5.60804786744919e-17 pua = -9.69608090826013e-25   ub = 1.57709603036933e-18 lub = 2.70418261178446e-25 wub = 1.90076613272594e-25 pub = -1.72042492405544e-31   uc = 5.27547128571428e-11 wuc = 2.5184628896543e-18   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0369023184564989 lu0 = 1.19547571570026e-09 wu0 = 7.85723699997298e-10 pu0 = 6.36693554141427e-16   a0 = -0.00563463721757884 la0 = 9.94339618217958e-07 wa0 = 1.67929185989264e-07 pa0 = -1.4805241581883e-13   keta = -0.0278164875170833 lketa = 1.51257770286112e-08 wketa = -5.3124783329442e-10 pketa = 4.68367214754356e-16   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 1.25311150817569e-07 lb0 = -3.98250176161571e-13 wb0 = -4.95051481262181e-14 pb0 = 1.14825829910165e-19   b1 = 8.91100461776685e-10 lb1 = -5.92828883505688e-15 wb1 = -2.67353263568358e-16 pb1 = 3.69016193641534e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.10519844832188+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.526923856721e-07 wnfactor = -2.29453106839087e-08 pnfactor = 1.09131759944877e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -1.51140947063948 lpclm = 2.61157244476481e-06 wpclm = 4.53904279422258e-07 ppclm = -4.86947979846725e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 4.02224876933938e-05 lalpha0 = 2.68300502765246e-12 walpha0 = -7.2082866296994e-12 palpha0 = -1.59090929518675e-18   alpha1 = 0.0   beta0 = 27.2922905296395 lbeta0 = 1.01342025956629e-05 wbeta0 = 1.05370642197692e-07 pbeta0 = -1.82069508834088e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37273   kt2 = -0.019151   at = 16473.456 lat = 0.006635672145984   ute = -1.0541754836 lute = -2.1549345294083e-7   ua1 = 3.0044e-9   ub1 = -4.31261405638e-18 lub1 = 1.05393077259064e-24 wub1 = 1.75292174856572e-25 pub1 = -3.2983606672842e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.81e-6   sbref = 2.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.85 nmos  lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.728386735310573+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.34637397725906e-08 wvth0 = 5.2666566987169e-08 pvth0 = -3.45482241506488e-14   k1 = 0.88325   k2 = -0.0291383388359659 lk2 = -1.30517583977133e-09 wk2 = -1.46848169712783e-09 pk2 = 6.32695408531147e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8492.84885669965 lvsat = 0.0694082954635248 wvsat = 0.0197290054408478 pvsat = -7.31450138659439e-9   ua = -3.82861509306095e-10 lua = 1.32555524410682e-16 wua = 1.41000568114642e-16 pua = -7.58382160644819e-23   ub = 2.32549915259295e-18 lub = -3.89400873886296e-25 wub = -5.11369612996666e-25 pub = 4.46377752737581e-31   uc = -1.61173239026743e-12 luc = 4.79314153221459e-17 wuc = 2.86119224374906e-17 puc = -2.30049333019162e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.031197658179612 lu0 = 6.2249095835737e-09 wu0 = 6.46411785925799e-09 pu0 = -4.36958315885253e-15   a0 = 1.1222   keta = -0.0552845267402473 lketa = 3.93425892571647e-08 wketa = 1.39656026395743e-08 pketa = -1.23125780487437e-14   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = -1.55109836393686e-06 lb0 = 1.07973280278847e-12 wb0 = 3.55901545683794e-13 pb0 = -2.42595305993719e-19   b1 = -2.57133129416897e-08 lb1 = 1.75271197803216e-14 wb1 = 1.727226837268e-14 pb1 = -1.17733999244801e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {1.08633246128656+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.36059452326231e-07 wnfactor = 6.79952258746182e-08 pnfactor = 2.8955309055563e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.74921264142699 lpclm = -1.14474539162902e-06 wpclm = -5.04773914435707e-07 ppclm = 3.58257228273436e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = -4.89943192907334e-06 lalpha0 = 4.24641137559259e-11 walpha0 = 1.09986774528583e-11 palpha0 = -1.76428242810766e-17   alpha1 = 0.0   beta0 = 28.1195549230774 lbeta0 = 9.40485652488993e-06 wbeta0 = 1.37871928038354e-06 pbeta0 = -2.9433250883165e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37954636 lkt1 = 6.00954836496017e-9   kt2 = -0.019151   at = 6959.10000000001 lat = 0.0150238709124   ute = -1.47412127 lute = 1.54745870397719e-7   ua1 = 6.387700286e-09 lua1 = -2.9828393309479e-15   ub1 = -7.6023113521e-18 lub1 = 3.95424633760003e-24 wub1 = -8.76460874282859e-25 pub1 = 5.97427284502672e-31   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.41e-6   sbref = 2.41e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.86 nmos  lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.756193750881052+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.4509476907191e-08 wvth0 = 1.26948451550699e-08 pvth0 = -7.30205956790419e-15   k1 = 0.88325   k2 = -0.0365971414389356 lk2 = 3.77901253130643e-09 wk2 = 8.0368156371074e-09 pk2 = -1.52198768407301e-16   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 69074.5339826344 lvsat = 0.0281136379410231 wvsat = 0.0284812536712035 pvsat = -1.32803488613411e-8   ua = -1.72394537052128e-10 lua = -1.09063406886232e-17 wua = 2.11892918410241e-17 pua = 5.82946304956173e-24   ub = -4.66126847511975e-19 lub = 1.51347190632123e-24 wub = 1.02070245067838e-24 pub = -5.97937720457623e-31   uc = 4.42120303724952e-11 luc = 1.66962889675873e-17 wuc = 2.52806521868463e-18 puc = -5.22523720271817e-24   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0292486307377091 lu0 = 7.55343685296258e-09 wu0 = 2.34845418748989e-09 pu0 = -1.56419863628321e-15   a0 = 1.1222   keta = 0.00243335972285715 wketa = -4.09767167214593e-9   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.792823767524713+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.59933603451776e-08 wnfactor = 1.56615574706987e-07 pnfactor = -3.14515110411376e-14   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = 2.23205414222425 lpclm = -7.9223154086647e-07 wpclm = -6.68355065865011e-07 ppclm = 4.69760030009101e-13   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 0.0001232773886929 lalpha0 = -4.49058215455533e-11 walpha0 = -3.55018893897525e-11 palpha0 = 1.40536360992533e-17   alpha1 = 0.0   beta0 = 47.254789997453 lbeta0 = -3.63840857026717e-06 wbeta0 = -5.59031623259135e-06 pbeta0 = 1.80702040260565e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.37073   kt2 = -0.019151   at = 6363.10800000001 lat = 0.015430120515312   ute = -1.12187464 lute = -8.53581134889591e-8   ua1 = 2.0117e-9   ub1 = -1.8012e-18   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 2.02e-6   sbref = 2.01e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_g5v0d10v5__model.87 nmos  lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 5.9182e-8   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 5.3521e-8   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -4.1292e-9   dwb = -1.6944e-9   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.794   rnoib = 0.38   tnoia = 7.50e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.2296e-08+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.2296e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {0.867132710849061+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.10772799840389e-08 wvth0 = -3.11206077793727e-08 pvth0 = 1.3801039921629e-14   k1 = 0.88325   k2 = -0.0111901330587341 lk2 = -8.45791735690028e-09 wk2 = 1.20499206834576e-08 pk2 = -2.08505463051124e-15   k3 = -0.884   dvt0 = 0.0   dvt1 = 0.53   dvt2 = -0.19251   dvt0w = 0.16   dvt1w = 6909100.0   dvt2w = -0.036016   w0 = 0.0   k3b = 0.43   phin = 0.0   lpe0 = 2.5e-8   lpeb = -2.182e-7   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 89887.224789178 lvsat = 0.0180894967917226 wvsat = 0.00811560157989138 pvsat = -3.47151765068993e-9   ua = -4.90459157183594e-10 lua = 1.42285030693016e-16 wua = 1.87364894706857e-16 pua = -7.42066896123266e-23   ub = 1.1862145118082e-18 lub = 7.17644823383695e-25 wub = -8.6222695918267e-25 pub = 3.08948868790214e-31   uc = 2.34878447920744e-10 luc = -7.51355217146811e-17 wuc = -4.0076299830518e-17 puc = 1.52945587621196e-23   rdsw = 724.62   prwb = 0.05626   prwg = 0.048   wr = 1.0   u0 = 0.0516028475882495 lu0 = -3.21315873406428e-09 wu0 = -6.58950363692804e-09 pu0 = 2.74064361843815e-15   a0 = 1.1222   keta = 0.0524023340347802 lketa = -2.40668569116974e-08 wketa = -1.97358619348568e-08 pketa = 7.53191540537099e-15   a1 = 0.0   a2 = 0.65972622   ags = 0.16025   b0 = 3.2933e-8   b1 = 0.0   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.20613+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}   nfactor = {0.093070007057392+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.0103324183126e-07 wnfactor = 3.28638900714631e-07 pnfactor = -1.14304137686155e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -8.0e-4   cdsc = 0.0   cdscb = 0.0   cdscd = 0.0   eta0 = 0.032   etab = -0.01932   dsub = 0.504   voffl = -4.2579486e-7   minv = 0.0   pclm = -0.211996235328686 lpclm = 3.84911106776619e-07 wpclm = 3.73761037308915e-07 ppclm = -3.21606014591758e-14   pdiblc1 = 0.21098   pdiblc2 = 2.0e-4   pdiblcb = -0.26831   drout = 0.36075   pscbe1 = 937310000.0   pscbe2 = 1.68e-6   pvag = 1.99   delta = 0.0246   alpha0 = 8.94787882294012e-05 lalpha0 = -2.86271988127158e-11 walpha0 = -3.04535189886956e-11 palpha0 = 1.16221591727698e-17   alpha1 = 0.0   beta0 = 50.1593290494611 lbeta0 = -5.03733914112016e-06 wbeta0 = -8.85477146394717e-06 pbeta0 = 3.37929956241495e-12   fprout = 10.125   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 5.06e-11   bgidl = 1058000000.0   cgidl = 4000.0   egidl = 0.8   aigbacc = 1.0   bigbacc = 0.0   cigbacc = 0.0   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = -0.383073607524285 lkt1 = 5.94512575356701e-09 wkt1 = -3.79395830272147e-08 pkt1 = 1.82730690108955e-14   kt2 = -0.019151   at = 66001.9113672411 lat = -0.0132940741832725 wat = -0.022015075377925 pat = 1.06032528447223e-8   ute = -2.56017331518108 lute = 6.07378307230558e-07 wute = 3.94065802376002e-07 pute = -1.89796276793168e-13   ua1 = -1.776800572e-09 lua1 = 1.82467826149579e-15   ub1 = -8.52358137256148e-18 lub1 = 3.23774087475502e-24 wub1 = 4.43437846422084e-24 pub1 = -2.13575630599347e-30   uc1 = -5.9821e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.6e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 0.89   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.0773   jss = 0.000375   jsws = 5.84e-11   xtis = 0.76   bvs = 12.636   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001344   tpbsw = 0.00099005   tpbswg = 0.0   tcj = 0.00067434   tcjsw = 0.0002493   tcjswg = 0.0   cgdo = 3.19377688e-10   cgso = 3.19377688e-10   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = 5.206e-11   cgdl = 5.206e-11   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = 4.867e-8   dwc = 3.2175e-8   vfbcv = -1.0   acde = 0.4176   moin = 15.0   noff = 4.0   voffcv = -0.4104   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.00099811712   mjs = 0.295   pbs = 0.72468   cjsws = 1.06590204e-10   mjsws = 0.037586   pbsws = 0.29067   cjswgs = 6.7554e-11   mjswgs = 0.78692   pbswgs = 0.54958   saref = 1.81e-6   sbref = 1.81e-6   wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__nfet_g5v0d10v5





















