** Translated using xdm 2.6.0 on Nov_14_2022_16_05_07_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* statistics {
* 	mismatch {
*     	}
*         process {
* 		vary sky130_fd_pr__res_xhigh_po__var_mult dist=gauss std=0.025
* 		vary sky130_fd_pr__res_high_po__var       dist=gauss std=0.025
*         }
* }
.SUBCKT sky130_fd_pr__res_xhigh_po r0 r1 sub PARAMS: W=1 L=1
* .param  mult = 1.0  rsheet = 2000.0   rend_mm = {0.0472/sqrt(w)}   leff = {l-0.0592}   weff = {w-0.056}   bp2 = -0.1228   bq2 = 1.304   bp22 = -0.2874   bp23 = 0.5252   sub1 = 1.2   sub2 = 41.26e-3   sub3 = 8.697e-3   sub4 = 24.0   sub5 = 39.86   body_pelgrom = 0.0347   res_match = {(body_pelgrom/sqrt(w*l*mult))*sky130_fd_pr__res_high_po__slope_spectre}   rhead0 = {188.2/(weff-0.0672*max(0.69-w,0)+1.41)}   rbody0 = {rsheet*leff/(weff-0.0672*max(0.69-w,0))}   rhead = {rhead0*(1+sky130_fd_pr__res_xhigh_po__var_mult)*(1+rend_mm/sqrt(mult)*sky130_fd_pr__res_high_po__con_slope_spectre)}   rbody = {rbody0*(1+sky130_fd_pr__res_xhigh_po__var_mult)*(1+res_match)}   Efac = {1/leff*(1+bp22/w+bp23*min(0.2,leff-0.5)*log(leff/w))}; HSpice Parser Retained (as a comment). Continuing.

* ;  Resistor voltco fitting parameters




* ;  Substrate voltco fitting parameters




* rend1 r0 t1 reshead r = {rhead}  tc1 = -4.3e-4   tc2 = -1.3e-5; HSpice Parser Retained (as a comment). Continuing.












*+ tnom = 25.0


* rend2 t2 r1 reshead r = {rhead}  tc1 = -4.3e-4   tc2 = -1.3e-5; HSpice Parser Retained (as a comment). Continuing.
*+ tnom = 25.0


* xc0 r0 r1 sub sky130_fd_pr__model__parasitic__res_po w = {w} l = {l}; HSpice Parser Retained (as a comment). Continuing.
* rbody t1 t2 r = {rbody*(1-bp2+bp2*sqrt(1+(bq2*abs(v(t1,t2))*Efac)**2))*  (sub1+sub2*tanh(sub3*(min(v(r0,sub)+v(r1,sub),sub4)+sub5))) / (sub1+sub2*tanh(sub3*sub5)) }   tc1 = -1.47e-3   tc2 = 2.7e-6; HSpice Parser Retained (as a comment). Continuing.
*+ tnom = 25.0



* .model resbody r tc1 = {-1.47e-3-5e-7*sky130_fd_pr__res_xhigh_po__var_mult*rsheet} tc2 = 2.7e-6 tnom = 25.0; HSpice Parser Retained (as a comment). Continuing.
.MODEL reshead R TC1=-4.3e-4 TC2=-1.3e-5 TNOM=25.0 LEVEL=1
.ENDS sky130_fd_pr__res_xhigh_po
