** Translated using xdm 2.6.0 on Nov_14_2022_16_05_05_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TOXE_MULT=1.042 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RSHP_MULT=1.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__OVERLAP_MULT=1.1981e+0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AJUNCTION_MULT=1.0559e+0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PJUNCTION_MULT=1.0542e+0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__WINT_DIFF=2.252e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__DLC_DIFF=-1.21275e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__DWC_DIFF=2.252e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_0=0.0066792 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_0=0.0055732 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_0=57405.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_0=-0.039836 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_0=-0.84048 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_0=1.8175e-9 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_0=-4.3477e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_0=-0.032489 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_1=0.11937 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_1=0.013842 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_1=-0.0048548 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_1=11004.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_1=0.050578 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_1=9.3332e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_1=0.59173 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_1=-2.2152e-18 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_2=5.2299e-2 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_2=9.1344e-3 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_2=-4.0166e-4 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_2=-1.2687e-2 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_2=2.4782e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_2=3.6143e+4 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_2=4.0028e-1 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_2=1.3690e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_3=2.0000e-2 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_3=6.1506e-3 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_3=5.9152e-3 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_3=-4.2250e-2 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_3=1.8174e-9 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_3=2.3364e+4 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_3=4.0000e-6 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_3=-5.2157e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_4=-0.049006 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_4=0.0067633 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_4=0.0052948 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_4=-0.042196 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_4=1.782e-9 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_4=47926.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_4=-1.0053 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_4=-4.6278e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_5=0.13767 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_5=0.014733 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_5=-0.0063472 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_5=0.06743 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_5=-2.5905e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_5=15839.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_5=0.62815 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_5=-2.734e-18 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_6=-2.9719e-18 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_6=0.15175 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_6=0.014735 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_6=-0.0073782 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_6=0.086313 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_6=-6.8974e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_6=27158.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_6=0.57872 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_7=-1.8438e-18 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_7=0.10854 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_7=0.013897 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_7=-0.0041489 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_7=0.035699 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_7=1.8882e-10 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_7=12478.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_7=0.60147 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_7=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
*




* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
.INCLUDE sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice























