** Translated using xdm 2.6.0 on Nov_14_2022_16_05_33_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 18
.PARAM 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__TOXE_MULT=0.948 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RBPB_MULT=0.8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__OVERLAP_MULT=8.6067e-1 SKY130_FD_PR__RF_NFET_01V8_LVT_B__AJUNCTION_MULT=8.2447e-1 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__PJUNCTION_MULT=7.5000e-1 SKY130_FD_PR__RF_NFET_01V8_LVT_B__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__RSHG_DIFF=-7.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__DLC_DIFF=1.1336e-8 SKY130_FD_PR__RF_NFET_01V8_LVT_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_B__XGW_DIFF=-6.4250e-8 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT_P42=0.85 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT_P42=0.65 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT_P42=0.65 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_CAP_MULT=0.85 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_DIST_MULT=0.75 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RGATE_STUB_MULT=0.75 SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RD_MULT=1.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT__AW_RS_MULT=1.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_0=-0.065542 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_0=0.0010442 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_0=-32505.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_0=-0.0038838 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_1=0.0043607 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_1=-0.059034 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_1=0.00085042 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_1=-26494.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_2=-0.0034116 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_2=-0.042789 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_2=0.0016287 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_2=-20516.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_3=0.016626 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_3=-0.073889 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_3=-0.0038 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_3=-37673.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_4=0.010615 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_4=-0.067217 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_4=-0.0036293 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_4=-25995.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_5=0.0050505 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_5=-0.029865 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_5=-0.00025925 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_5=-18682.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_6=0.0032612 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_6=-0.064411 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_6=-0.0093565 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_6=-31246.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_7=0.0089861 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_7=-0.056878 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_7=-0.0052178 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_7=-22366.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__UA_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__A0_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__NFACTOR_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__K2_DIFF_8=0.0046298 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VTH0_DIFF_8=-0.02487 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__U0_DIFF_8=-0.00059818 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__VSAT_DIFF_8=-16469.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM02__B1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_0=-0.0043971 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_0=-0.068994 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_0=-0.0051783 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_0=-28908.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_1=0.0032931 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_1=-0.066959 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_1=-0.0030718 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_1=-26301.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_2=0.0033757 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_2=-0.048089 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_2=-0.00068406 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_2=-15222.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_3=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_3=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_3=0.014866 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_3=-0.072281 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_3=-0.0047778 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_3=-38008.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_4=-0.008134 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_4=-24439.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_4=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_4=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_4=0.0080453 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_4=-0.062068 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_5=-0.041218 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_5=-0.0034389 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_5=-9878.8 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_5=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_5=0.0034441 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_6=0.0075537 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_6=-0.069722 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_6=-0.0070527 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_6=-35711.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_6=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_6=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_7=0.0046426 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_7=-0.055588 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_7=-0.0090538 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_7=-24756.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_7=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__PCLM_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__NFACTOR_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__A0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B0_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__K2_DIFF_8=0.0027331 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__U0_DIFF_8=-0.005212 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VSAT_DIFF_8=-7446.5 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__VTH0_DIFF_8=-0.041012 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__KT1_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__B1_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__AGS_DIFF_8=0.0 SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UB_DIFF_8=0.0 
+ SKY130_FD_PR__RF_NFET_01V8_LVT_BM04__UA_DIFF_8=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
*









* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
*















* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice















