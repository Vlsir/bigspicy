** Translated using xdm 2.6.0 on Nov_14_2022_16_05_31_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__NFET_05V0_NVT__TOXE_MULT=0.948 SKY130_FD_PR__NFET_05V0_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_05V0_NVT__OVERLAP_MULT=4.0927e-1 SKY130_FD_PR__NFET_05V0_NVT__AJUNCTION_MULT=5.6418e-1 
+ SKY130_FD_PR__NFET_05V0_NVT__PJUNCTION_MULT=8.4099e-1 SKY130_FD_PR__NFET_05V0_NVT__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__NFET_05V0_NVT__DLC_DIFF=3.0000e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__DWC_DIFF=-3.2175e-8 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_0=0.084235 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_0=-0.088752 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_0=-0.00071772 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_0=-0.010239 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_0=-3.0465e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_0=-0.042356 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_0=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_0=-0.0089574 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_0=-1.6353e-18 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_1=-1.3876e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_1=-0.036725 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_1=-0.051834 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_1=-0.0056229 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_1=-0.0086911 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_1=-2.5597e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_1=-0.025235 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_1=-0.0075728 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_2=-1.9312e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_2=0.12544 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_2=0.00061719 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_2=-0.011151 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_2=-4.1518e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_2=-7949.5 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_2=-0.043464 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_2=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_3=-1.9154e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_3=-0.0071658 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_3=-1.1337e-18 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_3=0.010177 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_3=0.0013249 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_3=-0.0054271 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_3=-0.0080273 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_3=-0.029234 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_4=-0.010027 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_4=-0.026425 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_4=-2.2287e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_4=-0.068222 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_4=-1.4787e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_4=-0.079945 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_4=-0.33061 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_4=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_4=-0.0024831 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_5=-0.0012384 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_5=-0.009243 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_5=-0.023314 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_5=-2.3342e-11 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_5=-0.017982 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_5=-1.3625e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_5=-0.012283 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_5=-0.089312 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_6=-0.072963 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_6=-0.0029725 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_6=-0.0083572 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_6=-0.029505 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_6=-2.0886e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_6=-0.013959 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_6=-1.2199e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_6=-0.042692 SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_7=0.079414 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_7=-8.6129e-5 
+ SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_7=-0.012564 SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_7=-0.049862 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_7=-3.2654e-11 
+ SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_7=-9440.5 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_7=-1.7558e-18 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_7=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_8=0.050854 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_8=2.7274e-7 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_8=-0.011083 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_8=-0.012082 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_8=-0.068342 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_8=-2.1309e-11 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_8=-2.2962e-8 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_8=-1.6897e-18 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_8=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_9=-0.15711 SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_9=-0.0083374 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_9=-0.012537 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_9=-0.057364 SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_9=-1.3616e-10 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_9=-13432.0 
+ SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_9=0.0 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_9=-1.1456e-18 SKY130_FD_PR__NFET_05V0_NVT__VSAT_DIFF_10=-11514.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VTH0_DIFF_10=-0.047797 SKY130_FD_PR__NFET_05V0_NVT__B0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KETA_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__B1_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__KT1_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__PCLM_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__NFACTOR_DIFF_10=0.058 
+ SKY130_FD_PR__NFET_05V0_NVT__AGS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__U0_DIFF_10=-0.012559 
+ SKY130_FD_PR__NFET_05V0_NVT__PDITS_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__K2_DIFF_10=0.0004686 
+ SKY130_FD_PR__NFET_05V0_NVT__UA_DIFF_10=-2.9266e-11 SKY130_FD_PR__NFET_05V0_NVT__ETA0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__UB_DIFF_10=-1.7087e-18 SKY130_FD_PR__NFET_05V0_NVT__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__VOFF_DIFF_10=0.0 SKY130_FD_PR__NFET_05V0_NVT__A0_DIFF_10=0.0 
+ SKY130_FD_PR__NFET_05V0_NVT__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0, L = 2.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0, L = 4.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0, L = 0.9
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0, L = 25.0
* -------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0, L = 2.0
* ------------------------------------
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0, L = 4.0
* ------------------------------------
*














* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0, L = 8.0
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0, L = 0.9
* ------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42, L = 1.0
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42, L = 0.9
* -------------------------------------
*




















* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7, L = 0.9
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_05v0_nvt.pm3.spice




















