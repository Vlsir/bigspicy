** Translated using xdm 2.6.0 on Nov_14_2022_16_05_26_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__res_iso_pw r0 r1 b
.PARAM 
+ L=-1 MULT=1.0 W=2.65 DL=0.52 AV=0.0133 BV=0.0302 TREF=30.0 LOCAL_VT=3.531e-3 UT=7.238e-6
Rpwres r0 r1 
+ R={rspwres*((l+dl)/w)*(1-av*(max(v(r0),v(r1))-min(v(r0),v(r1))))*(1+bv*(v(b)-min(v(r0),v(r1))))*(1+local_vt*(temp-tref)+ut*(temp-tref)*(temp-tref))}






.ENDS sky130_fd_pr__res_iso_pw

