** Translated using xdm 2.6.0 on Nov_14_2022_16_05_32_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 11
.PARAM 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TOXE_MULT=0.94 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RSHN_MULT=1.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__OVERLAP_MULT=0.76246 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AJUNCTION_MULT=8.1753e-1 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PJUNCTION_MULT=7.7786e-1 SKY130_FD_PR__ESD_NFET_G5V0D10V5__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__DLC_DIFF=1.7325e-8 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__DWC_DIFF=-3.2175e-8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_0=0.14328 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_0=-0.00045472 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_0=-0.0011699 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_0=-0.0040664 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_0=-7090.1 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_0=-8.363e-19 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_0=-2.0608e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_0=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_1=0.15647 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_1=0.00040364 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_1=0.00057999 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_1=-0.0025892 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_1=-6925.9 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_1=-7.4921e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_1=-1.8631e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_1=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_2=0.1669 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_2=2.8343e-5 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_2=-0.0010571 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_2=-0.0034839 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_2=-5424.6 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_2=-7.5872e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_2=1.2923e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_3=-1.6825e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_3=0.15401 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_3=0.0001604 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_3=-0.0013049 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_3=-0.0016799 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_3=-5330.1 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_3=-7.6166e-19 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_4=-8.2209e-19 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_4=-5.2787e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_4=0.14553 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_4=-0.0026632 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_4=-0.00096576 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_4=-0.0043485 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_4=-6212.8 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_5=-1.0249e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_5=1.3027e-10 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_5=0.17146 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_5=0.24441 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_5=-0.4 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_5=0.054151 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_5=-0.0059635 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_5=-3.7876e-5 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_6=-5.3272e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_6=-1.7366e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_6=0.14152 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_6=-0.0011048 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_6=-0.00069586 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_6=-0.0038289 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_6=-4075.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_7=-2741.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_7=-2.1212e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_7=2.6239e-12 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_7=0.12367 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_7=-0.0014188 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_7=-0.00098518 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_7=-0.0023054 SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_8=-0.0085839 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_8=-0.00047254 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_8=-1.1983e-18 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_8=1.2035e-10 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_8=0.17047 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_8=0.16645 SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_8=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_8=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_8=-0.39993 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_8=0.015735 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_9=-0.0059114 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_9=0.0013661 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_9=-0.010512 SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_9=-5727.6 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_9=7.8668e-20 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_9=-1.2856e-11 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_9=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_9=0.12716 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_9=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__KT1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__ETA0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UA_DIFF_10=6.7679e-12 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__BGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PCLM_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__CGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__TVOFF_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B1_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__AGIDL_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITSD_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VSAT_DIFF_10=-7615.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__UB_DIFF_10=-5.6629e-19 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__VOFF_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__B0_DIFF_10=0.0 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__K2_DIFF_10=-0.0031534 SKY130_FD_PR__ESD_NFET_G5V0D10V5__NFACTOR_DIFF_10=0.28192 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__A0_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__U0_DIFF_10=-0.00288 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__PDITS_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__VTH0_DIFF_10=-0.0017519 
+ SKY130_FD_PR__ESD_NFET_G5V0D10V5__KETA_DIFF_10=0.0 SKY130_FD_PR__ESD_NFET_G5V0D10V5__RDSW_DIFF_10=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
*
















* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
*























* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
.INCLUDE sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice























