** Translated using xdm 2.6.0 on Nov_14_2022_16_05_12_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* statistics {
*   mismatch {
*   }
* }
.SUBCKT sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4 c0 c1 b m4
* .param  mult = 1.0   ctot_a = {33.819e-15*sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor+0.0283/sqrt(6.8*6.1*mult*2)*33.819e-15*sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor*sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__slope}   cm4_c0 = {2.75e-15*c0m4m3_vpp}   cm4_c1 = {1.53e-15*c1m4m3_vpp}   cpl2s = {(6.51e-15-1.05e-15)*cpl2s_vpp}   rat_m3 = 0.12   rat_m2 = 0.37   rat_m1 = 0.37   rat_li = 0.12   rat_li2p = 0.02   cap_m3 = {rat_m3*ctot_a}   cap_m2 = {rat_m2*ctot_a}   cap_m1 = {rat_m1*ctot_a}   cap_li = {rat_li*ctot_a}   cap_li2p = {rat_li2p*ctot_a}   ll1 = 2.73   lm1 = 2.42   lm2 = 2.77   lm3 = 2.25   wl1 = 0.170   wm1 = 0.140   wm2 = 0.140   wm3 = 0.300   nfl1 = 34.0   nfm1 = 42.0   nfm2 = 38.0   nfm3 = 22.0   nvia2_c0 = 48.0   nvia2_c1 = 23.0   nvia_c0 = 60.0   nvia_c1 = 32.0   ncon_c0 = 64.0   ncon_c1 = 13.0   nlicon = 68.0; HSpice Parser Retained (as a comment). Continuing.

* ccmvpp6p8x6p1_polym4shield m4 b0  c = {cm4_c0}; HSpice Parser Retained (as a comment). Continuing.


































* cm4_1 m4 b1 c = {cm4_c1}; HSpice Parser Retained (as a comment). Continuing.
* rsm3 b0 b2 r = {rm3*lm3/wm3*(1/3)*(1/nfm3)}; HSpice Parser Retained (as a comment). Continuing.
* cm3 b2 b1 c = {cap_m3}; HSpice Parser Retained (as a comment). Continuing.
* rvia2_0 b0 c0 r = {rcvia2/nvia2_c0}; HSpice Parser Retained (as a comment). Continuing.
* rvia2_1 b1 c1 r = {rcvia2/nvia2_c1}; HSpice Parser Retained (as a comment). Continuing.
* rsm2 c0 c2 r = {rm2*lm2/wm2*(1/3)*(1/nfm2)}; HSpice Parser Retained (as a comment). Continuing.
* cm2 c2 c1 c = {cap_m2}; HSpice Parser Retained (as a comment). Continuing.
* rvia_0 c0 d0 r = {rcvia/nvia_c0}; HSpice Parser Retained (as a comment). Continuing.
* rvia_1 c1 d1 r = {rcvia/nvia_c1}; HSpice Parser Retained (as a comment). Continuing.
* rsm1 d0 d2 r = {rm1*lm1/wm1*(1/3)*(1/nfm1)}; HSpice Parser Retained (as a comment). Continuing.
* cm1 d2 d1 c = {cap_m1}; HSpice Parser Retained (as a comment). Continuing.
* rcon1 d0 e0 r = {rcl1/ncon_c0}; HSpice Parser Retained (as a comment). Continuing.
* rcon2 d1 e1 r = {rcl1/ncon_c1}; HSpice Parser Retained (as a comment). Continuing.
* rli1 e0 e2 r = {rl1*ll1/wl1*(1/3)*(1/nfl1)}; HSpice Parser Retained (as a comment). Continuing.
* cli e2 e1 c = {cap_li}; HSpice Parser Retained (as a comment). Continuing.
* rlicon e0 f0 r = {rcp1/nlicon}; HSpice Parser Retained (as a comment). Continuing.
* rpoly f0 f2 r = {rp1}; HSpice Parser Retained (as a comment). Continuing.
* cl12p e1 f2 c = {cap_li2p}; HSpice Parser Retained (as a comment). Continuing.
* cpl2b f0 b c = {cpl2s}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4
