** Translated using xdm 2.6.0 on Nov_14_2022_16_05_33_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_LVT__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__pfet_01v8_lvt d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.452509+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.64774   k2 = -0.04782713   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.0054e-9   ub = 3.0419e-18   uc = 4.9353e-11   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 0.0025322839   a0 = 1.75209   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 0.385036   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 0.0018466   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 0.01363   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60135   kt2 = -0.055045   at = 285600.0   ute = -0.22271   ua1 = 6.8217e-10   ub1 = -1.4864e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-0.452509+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.64774   k2 = -0.04782713   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.0054e-9   ub = 3.0419e-18   uc = 4.9353e-11   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 0.0025322839   a0 = 1.75209   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 0.385036   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 0.0018466   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 0.01363   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60135   kt2 = -0.055045   at = 285600.0   ute = -0.22271   ua1 = 6.8217e-10   ub1 = -1.4864e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.619357840e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.536148201e-8   k1 = 0.64774   k2 = -4.894119812e-02 lk2 = 8.906306163e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.064217540e-09 lua = 4.702109418e-16   ub = 3.130975120e-18 lub = -7.121021393e-25   uc = 3.779220780e-11 luc = 9.242159716e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.450704172e-03 lu0 = 6.521809796e-10   a0 = 1.841424756e+00 la0 = -7.141777734e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.685411252e-01 lags = 1.318666271e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 7.488388000e-05 lpdiblc2 = 1.416380735e-8   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 5.859893400e-03 ldelta = 6.211734020e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.113360000e-01 lkt1 = 7.983207840e-8   kt2 = -0.055045   at = 2.991709740e+05 lat = -1.084917945e-1   ute = -3.123143780e-01 lute = 7.163332395e-7   ua1 = 6.682694880e-10 lua1 = 1.111262531e-16   ub1 = -1.753625360e-19 lub1 = 2.136306418e-25   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.223840804e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.262384285e-8   k1 = 0.64774   k2 = -3.968662488e-02 lk2 = -2.806016118e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.566795664e+05 lvsat = -1.314939160e-1   ua = -3.113132120e-09 lua = 6.655953401e-16   ub = 3.175873360e-18 lub = -8.914436692e-25   uc = 6.136577640e-11 luc = -1.740665252e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.320245161e-03 lu0 = 1.173286451e-9   a0 = 2.262730999e+00 la0 = -2.397043431e-6   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.230875368e-01 lags = -8.601355939e-8   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.638259200e-04 lpdiblc2 = 1.340909727e-8   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.967986080e-02 ldelta = 6.914862420e-9   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.59135   kt2 = -0.055045   at = 3.780323040e+05 lat = -4.234954911e-1   ute = -0.13298   ua1 = 6.9609e-10   ub1 = -1.571260340e-19 lub1 = 1.407867582e-25   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos  lmin = 1.5e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.703903488e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.311985885e-8   k1 = 0.64774   k2 = -4.752564752e-02 lk2 = -1.242601443e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 90748.0   ua = -2.234840640e-09 lua = -1.086069188e-15   ub = 1.831961120e-18 lub = 1.788854902e-24   uc = 2.748768160e-11 luc = 6.582580702e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 3.154886244e-03 lu0 = -4.913217254e-10   a0 = 1.100574118e+00 la0 = -7.923774814e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.672471040e-01 lags = 4.242345998e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -3.278730240e-03 lpdiblc2 = 2.047437127e-8   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.696915040e-02 ldelta = 1.232110324e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.59135   kt2 = -0.055045   at = 2.058295840e+05 lat = -8.005438633e-2   ute = -0.13298   ua1 = 8.001002400e-10 lua1 = -2.074380227e-16   ub1 = -3.124733360e-19 lub1 = 4.506114173e-25   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos  lmin = 1e-06 lmax = 1.5e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.490338288e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.879532464e-8   k1 = 0.64774   k2 = -5.110258288e-02 lk2 = -7.080642224e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 9.002606560e+04 lvsat = 1.078858767e-3   ua = -3.153121440e-09 lua = 2.862096399e-16   ub = 3.140969440e-18 lub = -1.673271311e-25   uc = 6.937218560e-11 luc = 3.233604239e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.029192874e-03 lu0 = 1.190914448e-9   a0 = 8.695573776e-01 la0 = 2.659936693e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = -2.128955200e-02 lags = 7.059837785e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-1.529629600e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.324351258e-8   nfactor = {2.597759520e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.035070669e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 5.973280000e-04 lpdiblc2 = 1.468198984e-8   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.023634720e-02 ldelta = 2.238260434e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.510140000e-01 lkt1 = 8.916188160e-8   kt2 = -9.336122080e-02 lkt2 = 5.725976036e-8   at = 2.043466720e+05 lat = -7.783832264e-2   ute = 5.615488000e-02 lute = -2.826431647e-7   ua1 = 6.6129e-10   ub1 = -1.050445280e-20 lub1 = -6.508817357e-28   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.731173008e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.153279916e-9   k1 = 0.64774   k2 = -6.360790704e-02 lk2 = 5.354652121e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.327331360e+04 lvsat = 2.768179536e-2   ua = -2.789854560e-09 lua = -7.502294554e-17   ub = 2.825072160e-18 lub = 1.468011241e-25   uc = 7.576047360e-11 luc = -3.118909348e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 3.243992422e-03 lu0 = -1.708222323e-11   a0 = 1.205606459e+00 la0 = -6.817353743e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 9.534706400e-01 lags = -2.633177564e-7   b0 = 7.305551040e-07 lb0 = -7.264639954e-13   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.108370400e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.430647258e-8   nfactor = {2.476840480e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.989118669e-8   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -2.274734080e-02 lpdiblc2 = 3.789592849e-08 ppdiblc2 = 2.524354897e-29   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.136885600e-02 ldelta = 1.131243759e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -4.915308320e-01 lkt1 = -6.942818066e-8   kt2 = -1.576964320e-02 lkt2 = -1.989730440e-8   at = 1.920565792e+05 lat = -6.561705436e-2   ute = -5.958848000e-02 lute = -1.675479675e-7   ua1 = 4.288626720e-10 lua1 = 2.311257350e-16   ub1 = 5.703157168e-19 lub1 = -5.782184584e-25 wub1 = 2.295887404e-40 pub1 = 2.299005293e-46   uc1 = -2.284941472e-11 luc1 = 1.281623960e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos  lmin = 3.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.792412720e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 8.180971277e-9   k1 = 0.64774   k2 = -6.623966640e-02 lk2 = 6.655793948e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.582753360e+05 lvsat = -1.928720452e-2   ua = -3.074079200e-09 lua = 6.549771648e-17   ub = 3.030160000e-18 lub = 4.540569600e-26   uc = 8.394894400e-11 luc = -7.167289114e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.404704480e-03 lu0 = 3.978617355e-10   a0 = 1.223188640e+00 la0 = -7.686616762e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.111120000e-01 lags = 4.824355200e-9   b0 = -2.435183680e-06 lb0 = 8.386772594e-13   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -8.848803200e-02 lpdiblc2 = 7.039812622e-8   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.489701600e-02 ldelta = 9.568115290e-9   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.549200000e-01 lkt1 = 1.135142400e-8   kt2 = -0.056015   at = 1.376778160e+05 lat = -3.873219383e-2   ute = -0.39848   ua1 = 8.9635e-10   ub1 = -5.9922e-19   uc1 = 3.0734e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.44e-6   sbref = 1.44e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.865294601e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.376345466e-7   k1 = 0.64774   k2 = -5.280901249e-02 wk2 = 3.479868835e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.121800871e-09 wua = 8.130656698e-16   ub = 3.232079581e-18 wub = -1.328413503e-24   uc = 5.087094712e-11 wuc = -1.060293347e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.602789677e-03 wu0 = -4.924862376e-10   a0 = 1.746656298e+00 wa0 = 3.795467152e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.370225731e-01 wags = -3.631287082e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.350837605e-03 wpdiblc2 = -3.522123876e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 3.485427320e-03 wdelta = 7.086032711e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60135   kt2 = -0.055045   at = 285600.0   ute = -0.22271   ua1 = 6.8217e-10   ub1 = -1.4864e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.865294601e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.376345466e-7   k1 = 0.64774   k2 = -5.280901249e-02 wk2 = 3.479868835e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.121800871e-09 wua = 8.130656698e-16   ub = 3.232079581e-18 wub = -1.328413503e-24   uc = 5.087094712e-11 wuc = -1.060293347e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.602789677e-03 wu0 = -4.924862376e-10   a0 = 1.746656298e+00 wa0 = 3.795467152e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.370225731e-01 wags = -3.631287082e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.350837605e-03 wpdiblc2 = -3.522123876e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 3.485427320e-03 wdelta = 7.086032711e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60135   kt2 = -0.055045   at = 285600.0   ute = -0.22271   ua1 = 6.8217e-10   ub1 = -1.4864e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.981316602e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.275262867e-08 wvth0 = 2.528299327e-07 pvth0 = -1.214779942e-13   k1 = 0.64774   k2 = -5.805719263e-02 lk2 = 4.195605127e-08 wk2 = 6.367565923e-08 pk2 = -2.308540559e-13   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.327222541e-09 lua = 1.642222999e-15 wua = 1.837102555e-15 pua = -8.186560478e-21   ub = 3.543176576e-18 lub = -2.487033812e-24 wub = -2.879246953e-24 pub = 1.239798293e-29   uc = 1.049460290e-11 luc = 3.227846462e-16 wuc = 1.906750805e-16 puc = -1.609096955e-21   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.370302029e-03 lu0 = 1.858599252e-09 wu0 = 5.616128242e-10 pu0 = -8.426889539e-15   a0 = 2.069238474e+00 la0 = -2.578850947e-06 wa0 = -1.591289752e-06 pa0 = 1.302483162e-11   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.890458391e-01 lags = -4.158947976e-07 wags = -8.417312105e-07 pags = 3.826139844e-12   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.270175929e-04 lpdiblc2 = 1.980896560e-08 wpdiblc2 = 1.410291480e-09 ppdiblc2 = -3.943170132e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -1.193099316e-02 ldelta = 1.232450319e-07 wdelta = 1.242701966e-07 pdelta = -4.269798606e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.113360000e-01 lkt1 = 7.983207840e-8   kt2 = -0.055045   at = 2.991709740e+05 lat = -1.084917945e-1   ute = -3.123143780e-01 lute = 7.163332395e-7   ua1 = 6.682694880e-10 lua1 = 1.111262531e-16   ub1 = -1.753625360e-19 lub1 = 2.136306418e-25   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.970759399e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.109043407e-07 wvth0 = -1.767785765e-07 pvth0 = 1.594550235e-12   k1 = 0.64774   k2 = -2.489203631e-02 lk2 = -9.051884911e-08 wk2 = -1.033409113e-07 pk2 = 4.362769332e-13   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 2.387323757e+05 lvsat = -4.592456576e-01 wvsat = -5.731428116e-01 pvsat = 2.289361647e-6   ua = -3.645202145e-09 lua = 2.912360732e-15 wua = 3.716534667e-15 pua = -1.569376411e-20   ub = 3.994770385e-18 lub = -4.290880126e-24 wub = -5.720035029e-24 pub = 2.374522682e-29   uc = 1.110001615e-10 luc = -7.867475726e-17 wuc = -3.466985627e-16 puc = 5.373883255e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.830227593e-03 lu0 = 4.015872580e-09 wu0 = 3.422796234e-09 pu0 = -1.985560055e-14   a0 = 3.513946251e+00 la0 = -8.349591691e-06 wa0 = -8.739798589e-06 pa0 = 4.157883532e-11   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 6.916239938e-01 lags = -1.225072979e-06 wags = -1.875740042e-06 pags = 7.956384720e-12   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.375208404e-03 lpdiblc2 = 9.814074073e-09 wpdiblc2 = -1.474810800e-08 ppdiblc2 = 2.511140956e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 3.346518452e-02 ldelta = -5.808546025e-08 wdelta = -9.629114790e-08 pdelta = 4.540303739e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.59135   kt2 = -0.055045   at = 5.814493013e+05 lat = -1.236024345e+00 wat = -1.420877490e+00 pat = 5.675553047e-6   ute = -0.13298   ua1 = 6.9609e-10   ub1 = -2.449776196e-19 lub1 = 4.917011319e-25 wub1 = 6.136475426e-25 pub1 = -2.451153744e-30   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos  lmin = 1.5e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-6.295995097e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.528406671e-07 wvth0 = 1.112083631e-06 pvth0 = -9.759565522e-13   k1 = 0.64774   k2 = -5.921996873e-02 lk2 = -2.205522070e-08 wk2 = 8.168539499e-08 pk2 = 6.726046804e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -3.876929948e+05 lvsat = 7.900971013e-01 wvsat = 3.341933314e+00 pvsat = -5.518866177e-6   ua = -4.901468211e-10 lua = -3.380081607e-15 wua = -1.218677007e-14 pua = 1.602378686e-20   ub = -8.162212032e-19 lub = 5.304161498e-24 wub = 1.849768064e-23 pub = -2.455458531e-29   uc = 5.303659099e-11 luc = 3.692778787e-17 wuc = -1.784603584e-16 puc = 2.018540508e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 5.342101450e-03 lu0 = -2.988208640e-09 wu0 = -1.527780319e-08 pu0 = 1.744087495e-14   a0 = -7.730963958e-01 la0 = 2.004861626e-07 wa0 = 1.308767848e-05 pa0 = -1.953884943e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.710450387e-01 lags = -5.857103109e-07 wags = -1.423538356e-06 pags = 7.054513679e-12   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -6.755076593e-03 lpdiblc2 = 2.802351447e-08 wpdiblc2 = 2.428244614e-08 ppdiblc2 = -5.273112762e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -6.396132487e-03 ldelta = 2.141395040e-08 wdelta = 1.632076225e-07 pdelta = -6.351397383e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -8.148396719e-01 lkt1 = 4.457278017e-07 wkt1 = 1.561086086e-06 pkt1 = -3.113430090e-12   kt2 = -2.067721383e-01 lkt2 = 3.026046046e-07 wkt2 = 1.059821344e-06 pkt2 = -2.113707688e-12   at = -8.460038989e+05 lat = 1.610888317e+00 wat = 7.347107366e+00 pat = -1.181131595e-5   ute = -0.13298   ua1 = 8.464370986e-10 lua1 = -2.998522535e-16 wua1 = -3.236651818e-16 pua1 = 6.455178386e-22   ub1 = 3.893300660e-20 lub1 = -7.453022106e-26 wub1 = -2.454590171e-24 pub1 = 3.668139551e-30   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos  lmin = 1e-06 lmax = 1.5e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.992457806e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.195994570e-08 wvth0 = 3.507328936e-07 pvth0 = 1.618059900e-13   k1 = 0.64774   k2 = -5.528005725e-02 lk2 = -2.794302442e-08 wk2 = 2.917985900e-08 pk2 = 1.457247410e-13   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 4.247553090e+05 lvsat = -4.240256438e-01 wvsat = -2.338099832e+00 pvsat = 2.969375355e-6   ua = -3.222586688e-09 lua = 7.032765301e-16 wua = 4.852180921e-16 pua = -2.913232247e-21   ub = 3.124193358e-18 lub = -5.843940213e-25 wub = 1.171817404e-25 pub = 2.913232247e-30   uc = 1.040374915e-10 luc = -3.928795792e-17 wuc = -2.421388260e-16 puc = 2.970151527e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.765272969e-03 lu0 = 2.357003841e-09 wu0 = 1.843493200e-09 pu0 = -8.145190384e-15   a0 = -2.280614091e+00 la0 = 2.453320606e-06 wa0 = 2.200409891e-05 pa0 = -1.527858364e-11   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = -1.808012019e+00 lags = 2.670672557e-06 wags = 1.248034220e-05 pags = -1.372344542e-11   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-8.083669331e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.510290055e-07 wvoff = -5.038054349e-07 pvoff = 7.528868419e-13   nfactor = {2.748456325e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.155520115e-07 wnfactor = -1.052624414e-06 pnfactor = 1.573041924e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 1.739099758e-02 lpdiblc2 = -8.060378777e-09 wpdiblc2 = -1.173045881e-07 ppdiblc2 = 1.588565364e-13   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 5.502178720e-03 ldelta = 3.633114129e-09 wdelta = 3.306839408e-08 pdelta = 1.309660891e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.258095973e-01 lkt1 = 1.632412582e-07 wkt1 = -1.760539626e-07 pkt1 = -5.174480013e-13   kt2 = 5.836591748e-02 lkt2 = -9.361770594e-08 wkt2 = -1.059821344e-06 pkt2 = 1.053886344e-12   at = 9.371843412e+05 lat = -1.053908189e+00 wat = -5.118906295e+00 pat = 6.817894865e-6   ute = 3.430240933e-01 lute = -7.113405170e-07 wute = -2.003795225e-06 pute = 2.994471584e-12   ua1 = 5.166036478e-10 lua1 = 1.930508554e-16 wua1 = 1.010641115e-15 pua1 = -1.348469491e-21   ub1 = -9.418840951e-21 lub1 = -2.273220083e-27 wub1 = -7.583050876e-27 pub1 = 1.133211123e-32   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-5.702377328e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.863445151e-08 wvth0 = 6.783908790e-07 pvth0 = -1.640171107e-13   k1 = 0.64774   k2 = -1.117953342e-01 lk2 = 2.825576697e-08 wk2 = 3.365914916e-07 pk2 = -1.599653865e-13   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 8.779420910e+03 lvsat = -1.037922070e-02 wvsat = 3.806424561e-01 pvsat = 2.658580241e-7   ua = -1.775445946e-09 lua = -7.357602237e-16 wua = -7.085692860e-15 pua = 4.615281603e-21   ub = 1.488559256e-18 lub = 1.042080530e-24 wub = 9.335606789e-24 pub = -6.253569621e-30   uc = 3.651704314e-11 luc = 2.785437597e-17 wuc = 2.741172454e-16 puc = -2.163498847e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 5.222720488e-03 lu0 = -1.081081971e-09 wu0 = -1.382151052e-08 pu0 = 7.432089310e-15   a0 = 8.974429753e-01 la0 = -7.069393404e-07 wa0 = 2.152536727e-06 pa0 = 4.461809795e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.132073412e+00 lags = -2.529483965e-07 wags = -1.247548938e-06 pags = -7.243047650e-14   b0 = -5.063575781e-07 lb0 = 5.035219756e-13 wb0 = 8.639894456e-12 pb0 = -8.591511047e-18   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-2.829633067e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.996569883e-08 wvoff = 5.038054349e-07 pvoff = -2.490814070e-13   nfactor = {2.326143675e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.043956869e-07 wnfactor = 1.052624414e-06 pnfactor = -5.204175102e-13   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -4.153656099e-02 lpdiblc2 = 5.053718547e-08 wpdiblc2 = 1.312436049e-07 ppdiblc2 = -8.829978676e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 4.106256910e-03 ldelta = 5.021218777e-09 wdelta = 1.205800832e-07 pdelta = 4.394446541e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -3.088218836e-01 lkt1 = -1.519713243e-07 wkt1 = -1.276230775e-06 pkt1 = 5.765678205e-13   kt2 = -1.576964320e-02 lkt2 = -1.989730440e-8   at = -3.026155963e+05 lat = 1.789488692e-01 wat = 3.455308890e+00 pat = -1.708304715e-6   ute = -3.464576933e-01 lute = -2.571982844e-08 wute = 2.003795225e-06 pute = -9.906763590e-13   ua1 = 5.272121655e-10 lua1 = 1.825017454e-16 wua1 = -6.869759332e-16 pua1 = 3.396409014e-22   ub1 = 5.692301050e-19 lub1 = -5.776817319e-25 wub1 = 7.583050876e-27 pub1 = -3.749060353e-33   uc1 = -2.284941472e-11 luc1 = 1.281623960e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos  lmin = 3.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-5.648983947e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.599468275e-08 wvth0 = 5.983191133e-07 pvth0 = -1.244296297e-13   k1 = 0.64774   k2 = -6.003801544e-02 lk2 = 2.666948580e-09 wk2 = -4.331882962e-08 pk2 = 2.786227636e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.612834642e+05 lvsat = 1.231398697e-01 wvsat = 2.930638358e+00 pvsat = -9.948599499e-7   ua = -4.135503596e-09 lua = 4.310522785e-16 wua = 7.414100356e-15 pua = -2.553416163e-21   ub = 4.593542837e-18 lub = -4.930233532e-25 wub = -1.092030416e-23 pub = 3.760952753e-30   uc = 1.610911660e-10 luc = -3.373507037e-17 wuc = -5.388421234e-16 puc = 1.855772273e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.348473447e-03 lu0 = 8.343457659e-10 wu0 = 7.377824465e-09 pu0 = -3.048861904e-15   a0 = -4.050956890e+00 la0 = 1.739549553e-06 wa0 = 3.684015968e-05 pa0 = -1.268775100e-11   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.093466766e+00 lags = -2.338612706e-07 wags = -4.766280794e-06 pags = 1.667230553e-12   b0 = 1.687858594e-06 lb0 = -5.812984996e-13 wb0 = -2.879964819e-11 pb0 = 9.918598835e-18   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.576217744e-01 lpdiblc2 = 1.079297150e-07 wpdiblc2 = 4.829025089e-07 ppdiblc2 = -2.621599489e-13   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.427768939e-03 ldelta = 6.345463229e-09 wdelta = 1.639338172e-07 pdelta = 2.251037933e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.029989305e-01 lkt1 = -6.530192349e-09 wkt1 = -3.626711629e-07 pkt1 = 1.249039485e-13   kt2 = -0.056015   at = 1.376778160e+05 lat = -3.873219383e-2   ute = -0.39848   ua1 = 8.9635e-10   ub1 = -5.9922e-19   uc1 = 3.0734e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.44e-6   sbref = 1.44e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.449641247e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.042935440e-8   k1 = 0.64774   k2 = -4.424453353e-02 wk2 = -7.895650373e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.107952400e-09 wua = 7.440303781e-16   ub = 3.070076680e-18 wub = -5.208212647e-25   uc = 3.055610254e-11 wuc = 9.066754188e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.148846437e-03 wu0 = 1.770442606e-9   a0 = 1.766947499e+00 wa0 = -6.319794032e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.736102592e-01 wags = -4.701527959e-8   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 7.438602708e-04 wpdiblc2 = 4.488735271e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.327168129e-02 wdelta = 2.207538132e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60135   kt2 = -0.055045   at = 2.898686186e+05 wat = -2.127926881e-2   ute = -1.196661430e-01 wute = -5.136785731e-7   ua1 = 6.8217e-10   ub1 = -1.464161392e-19 wub1 = -1.108605263e-26   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.449641247e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.042935440e-8   k1 = 0.64774   k2 = -4.424453353e-02 wk2 = -7.895650373e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.107952400e-09 wua = 7.440303781e-16   ub = 3.070076680e-18 wub = -5.208212647e-25   uc = 3.055610254e-11 wuc = 9.066754188e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.148846437e-03 wu0 = 1.770442606e-9   a0 = 1.766947499e+00 wa0 = -6.319794032e-8   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.736102592e-01 wags = -4.701527959e-8   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 7.438602708e-04 wpdiblc2 = 4.488735271e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.327168129e-02 wdelta = 2.207538132e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.60135   kt2 = -0.055045   at = 2.898686186e+05 wat = -2.127926881e-2   ute = -1.196661430e-01 wute = -5.136785731e-7   ua1 = 6.8217e-10   ub1 = -1.464161392e-19 wub1 = -1.108605263e-26   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.387610425e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.958991985e-08 wvth0 = -4.313544628e-08 pvth0 = 5.881064426e-13   k1 = 0.64774   k2 = -3.687425423e-02 lk2 = -5.892096088e-08 wk2 = -4.192230550e-08 pk2 = 2.720226917e-13   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.152665434e-09 lua = 3.574538789e-16 wua = 9.669269988e-16 pua = -1.781924744e-21   ub = 3.070076680e-18 wub = -5.208212647e-25   uc = 3.055610254e-11 wuc = 9.066754188e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.895206273e-03 lu0 = 2.027700927e-09 wu0 = 2.929987976e-09 pu0 = -9.269869507e-15   a0 = 1.823456539e+00 la0 = -4.517558671e-07 wa0 = -3.660550087e-07 pa0 = 2.421160548e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.208830350e-01 lags = 4.215225210e-07 wags = -3.431560364e-09 pags = -3.484256850e-13   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.497520522e-03 lpdiblc2 = 1.791849461e-08 wpdiblc2 = 8.242314363e-09 ppdiblc2 = -3.000761269e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.181842103e-02 ldelta = 1.161794385e-08 wdelta = 5.878226883e-09 pdelta = 1.294865314e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.113360000e-01 lkt1 = 7.983207840e-8   kt2 = -0.055045   at = 3.077022352e+05 lat = -1.425690643e-01 wat = -4.252874665e-02 pat = 1.698768256e-7   ute = -1.063709255e-01 lute = -1.062872873e-07 wute = -1.026637996e-06 pute = 4.100802812e-12   ua1 = 6.682694880e-10 lua1 = 1.111262531e-16   ub1 = -1.709179279e-19 lub1 = 1.958770991e-25 wub1 = -2.215658479e-26 pub1 = 8.850226230e-32   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.472146933e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.582265732e-08 wvth0 = 7.316551589e-08 pvth0 = 1.235538793e-13   k1 = 0.64774   k2 = -5.566791247e-02 lk2 = 1.614842762e-08 wk2 = 5.007830862e-08 pk2 = -9.546456129e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.916032420e-09 lua = -5.877530322e-16 wua = 8.158858559e-17 pua = 1.754471013e-21   ub = 2.775291051e-18 lub = 1.177491717e-24 wub = 3.591279877e-25 pub = -3.514869294e-30   uc = -2.128076763e-12 luc = 1.305536858e-16 wuc = 2.172511354e-16 puc = -5.056255061e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.375100637e-03 lu0 = 1.108108785e-10 wu0 = 7.065779573e-10 pu0 = -3.886805294e-16   a0 = 1.388012170e+00 la0 = 1.287583117e-06 wa0 = 1.858084846e-06 pa0 = -6.462943686e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 2.179597572e-01 lags = 8.326392618e-07 wags = 4.854989135e-07 pags = -2.301409570e-12   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.467300553e-03 lpdiblc2 = 1.779778396e-08 wpdiblc2 = 4.406983594e-09 ppdiblc2 = -1.468776747e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.266017464e-02 ldelta = 8.255643234e-09 wdelta = 7.422825020e-09 pdelta = 1.233167886e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.59135   kt2 = -0.055045   at = 2.853630531e+05 lat = -5.333743550e-02 wat = 5.512666901e-02 pat = -2.201979667e-7   ute = -0.13298   ua1 = 6.9609e-10   ub1 = -1.2188e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos  lmin = 1.5e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.382725820e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.365680408e-08 wvth0 = 1.583097125e-07 pvth0 = -4.625770650e-14   k1 = 0.64774   k2 = -5.250534235e-02 lk2 = 9.840997767e-09 wk2 = 4.821266018e-08 pk2 = -9.174371205e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.199177925e+05 lvsat = -7.900971013e-01 wvsat = -1.182550026e+00 pvsat = 2.358477772e-6   ua = -3.003633671e-09 lua = -4.130410963e-16 wua = 3.430825262e-16 pua = 1.232947498e-21   ub = 2.892636887e-18 lub = 9.434571803e-25 wub = 8.845033135e-27 pub = -2.816264969e-30   uc = -3.342407414e-11 luc = 1.929704230e-16 wuc = 2.525502073e-16 puc = -5.760259751e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.919212887e-03 lu0 = 1.020033408e-09 wu0 = 1.785460591e-09 pu0 = -2.540404054e-15   a0 = 1.832594506e+00 la0 = 4.009081077e-07 wa0 = 9.818426055e-08 pa0 = -2.952997960e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = -1.301370049e-01 lags = 1.526883444e-06 wags = 1.074878188e-06 pags = -3.476867595e-12   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -7.423973215e-03 lpdiblc2 = 2.967777192e-08 wpdiblc2 = 2.761692791e-08 ppdiblc2 = -6.097768041e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -1.440346889e-02 ldelta = 6.223137389e-08 wdelta = 2.031245788e-07 pdelta = -2.669907892e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -3.678603281e-01 lkt1 = -4.457278017e-07 wkt1 = -6.671273982e-07 pkt1 = 1.330518883e-12   kt2 = 9.668213828e-02 lkt2 = -3.026046046e-07 wkt2 = -4.529127907e-07 pkt2 = 9.032892697e-13   at = 1.110114556e+06 lat = -1.698221833e+00 wat = -2.404237026e+00 pat = 4.684756987e-6   ute = -0.13298   ua1 = 9.090011608e-10 lua1 = -4.246300191e-16 wua1 = -6.355500347e-16 pua1 = 1.267540989e-21   ub1 = -9.483448068e-19 lub1 = 1.648301411e-24 wub1 = 2.467037119e-24 pub1 = -4.920258829e-30   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos  lmin = 1e-06 lmax = 1.5e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.838287605e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.442234913e-08 wvth0 = 2.738783084e-07 pvth0 = -2.189634161e-13   k1 = 0.64774   k2 = -3.886579843e-02 lk2 = -1.054193667e-08 wk2 = -5.264600912e-08 pk2 = 5.897948335e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -2.950518845e+05 lvsat = 4.277935839e-01 wvsat = 1.250173578e+00 pvsat = -1.276984382e-6   ua = -3.161590542e-09 lua = -1.769903496e-16 wua = 1.811493738e-16 pua = 1.474940401e-21   ub = 3.631122076e-18 lub = -1.601350853e-25 wub = -2.409882253e-24 pub = 7.982810867e-31   uc = 1.588360267e-10 luc = -9.434307180e-17 wuc = -5.153121542e-16 puc = 5.714675381e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 3.556774614e-03 lu0 = -1.427138838e-09 wu0 = -7.087228491e-09 pu0 = 1.071894251e-14   a0 = 2.670256879e+00 la0 = -8.508945424e-07 wa0 = -2.676230509e-06 pa0 = 1.193087472e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.218875403e+00 lags = -4.890806979e-07 wags = -2.608836892e-06 pags = 2.028076221e-12   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {6.773703047e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.330880713e-06 wnfactor = -2.111867254e-05 pnfactor = 3.155974424e-11   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.483574667e-02 lpdiblc2 = 4.075392618e-08 wpdiblc2 = 4.334727888e-08 ppdiblc2 = -8.448511689e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 3.774569402e-02 ldelta = -1.570033516e-08 wdelta = -1.276670774e-07 pdelta = 2.273442618e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -8.543183066e-01 lkt1 = 2.812350014e-07 wkt1 = 9.630729214e-07 pkt1 = -1.105652475e-12   kt2 = -2.450883591e-01 lkt2 = 2.081372267e-07 wkt2 = 4.529127907e-07 pkt2 = -4.503764790e-13   at = -6.458038851e+05 lat = 9.258226854e-01 wat = 2.772365996e+00 pat = -3.051158569e-6   ute = -6.691962966e-01 lute = 8.013216337e-07 wute = 3.042172006e-06 pute = -4.546221845e-12   ua1 = 5.918468712e-10 lua1 = 4.932535128e-17 wua1 = 6.355500347e-16 pua1 = -6.319909545e-22   ub1 = 4.839473348e-19 lub1 = -4.921159657e-25 wub1 = -2.467037119e-24 pub1 = 2.453221711e-30   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.211650916e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.789040322e-08 wvth0 = -6.474339260e-08 pvth0 = 1.177620033e-13   k1 = 0.64774   k2 = -4.217404180e-02 lk2 = -7.252219466e-09 wk2 = -1.047399277e-08 pk2 = 1.704363029e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.809084120e+04 lvsat = 1.164044575e-01 wvsat = 3.342245790e-01 pvsat = -3.661646974e-7   ua = -3.860260525e-09 lua = 5.177670821e-16 wua = 3.307207888e-15 pua = -1.633612185e-21   ub = 4.002440454e-18 lub = -5.293740804e-25 wub = -3.196211651e-24 pub = 1.580207040e-30   uc = 7.475688874e-11 luc = -1.073477697e-17 wuc = 8.348977963e-17 puc = -2.398110499e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 7.659748549e-04 lu0 = 1.348032443e-09 wu0 = 8.395580388e-09 pu0 = -4.677162639e-15   a0 = 1.714069737e+00 la0 = 9.993795093e-08 wa0 = -1.918386880e-06 pa0 = 4.394877672e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.057449275e+00 lags = -3.285585568e-07 wags = -8.755440330e-07 pags = 3.044898019e-13   b0 = 1.436664019e-06 lb0 = -1.428618701e-12 wb0 = -1.046161472e-12 pb0 = 1.040302968e-18   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {4.071697472e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.061880156e-5   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -9.804184284e-03 lpdiblc2 = 3.575054054e-08 wpdiblc2 = -2.694381612e-08 ppdiblc2 = -1.458765203e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.953963187e-03 ldelta = 1.889656198e-08 wdelta = 1.263243228e-07 pdelta = -2.522478645e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.349831360e-01 lkt1 = -3.631189225e-08 wkt1 = -1.488060756e-07 pkt1 = -1.615587134e-27   kt2 = -8.330096427e-03 lkt2 = -2.729518971e-08 wkt2 = -3.708649776e-08 pkt2 = 3.687881337e-14   at = 5.138530430e+05 lat = -2.273401638e-01 wat = -6.148264673e-01 pat = 3.170656163e-7   ute = 6.128402314e-01 lute = -4.735354898e-07 wute = -2.778350976e-06 pute = 1.241706208e-12   ua1 = 3.894048800e-10 lua1 = 2.506336673e-16   ub1 = 5.176959761e-19 lub1 = -5.256756146e-25 wub1 = 2.644831570e-25 pub1 = -2.630020513e-31   uc1 = -2.284941472e-11 luc1 = 1.281623960e-17 wuc1 = 2.465190329e-32 puc1 = 1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos  lmin = 3.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.077983629e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.449891392e-08 wvth0 = -1.848320861e-07 pvth0 = 1.771338534e-13   k1 = 0.64774   k2 = -5.005687440e-02 lk2 = -3.354947025e-09 wk2 = -9.307529680e-08 pk2 = 5.788171500e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 6.576482278e+05 lvsat = -1.997927144e-01 wvsat = -1.650280235e+00 pvsat = 6.149744828e-7   ua = -2.883571214e-09 lua = 3.489188677e-17 wua = 1.173157339e-15 pua = -5.785375939e-22   ub = 2.725739067e-18 lub = 1.018270854e-25 wub = -1.609212711e-24 pub = 7.955947642e-31   uc = -1.338483519e-11 luc = 3.284249134e-17 wuc = 3.309291173e-16 puc = -1.463151135e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.516996829e-03 lu0 = 4.823271788e-10 wu0 = 1.552679318e-09 pu0 = -1.294032350e-15   a0 = 5.712683402e+00 la0 = -1.876976645e-06 wa0 = -1.183205582e-05 pa0 = 5.340805693e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = -1.142113310e-01 lags = 2.507104469e-07 wags = 1.254052488e-06 pags = -7.483827182e-13   b0 = -4.788880065e-06 lb0 = 1.649290294e-12 wb0 = 3.487204908e-12 pb0 = -1.200993370e-18   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {4.071697472e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.061880156e-5   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -3.097773221e-02 lpdiblc2 = 4.621874263e-08 wpdiblc2 = -1.484241202e-07 ppdiblc2 = 4.547221030e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 5.923589745e-02 ldelta = -8.929226321e-09 wdelta = -1.242424782e-07 pdelta = 9.865543992e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.801685910e-01 lkt1 = 3.546779672e-08 wkt1 = 2.202329919e-08 pkt1 = -8.445804291e-14   kt2 = -8.081348924e-02 lkt2 = 8.540599695e-09 wkt2 = 1.236216592e-07 pkt2 = -4.257529943e-14   at = 1.201648976e+05 lat = -3.270074473e-02 wat = 8.730273890e-02 pat = -3.006706328e-8   ute = -2.220717825e-01 lute = -6.075499010e-08 wute = -8.794034317e-07 pute = 3.028665419e-13   ua1 = 8.9635e-10   ub1 = -4.223690402e-19 lub1 = -6.090747055e-26 wub1 = -8.816105234e-25 pub1 = 3.036266643e-31   uc1 = 3.0734e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.44e-6   sbref = 1.44e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.499316648e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.525770017e-8   k1 = 0.64774   k2 = -5.094469785e-02 wk2 = 1.210466172e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.845106338e-09 wua = -4.057773476e-17   ub = 2.873731934e-18 wub = 6.527722548e-26   uc = 5.912933226e-11 wuc = 5.375079648e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.832952674e-03 wu0 = -2.716473513e-10   a0 = 1.879412537e+00 wa0 = -3.989114773e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.985572581e-01 wags = -1.214832690e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.668905030e-03 wpdiblc2 = -1.257615736e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.448898624e-02 wdelta = -1.140881238e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.914995200e-01 wkt1 = -2.940415562e-8   kt2 = -0.055045   at = 2.869166035e+05 wat = -1.246736198e-2   ute = -0.29175   ua1 = 6.8217e-10   ub1 = -1.5013e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.499316648e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.525770017e-8   k1 = 0.64774   k2 = -5.094469785e-02 wk2 = 1.210466172e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.845106338e-09 wua = -4.057773476e-17   ub = 2.873731934e-18 wub = 6.527722548e-26   uc = 5.912933226e-11 wuc = 5.375079648e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.832952674e-03 wu0 = -2.716473513e-10   a0 = 1.879412537e+00 wa0 = -3.989114773e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.985572581e-01 wags = -1.214832690e-7   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.668905030e-03 wpdiblc2 = -1.257615736e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.448898624e-02 wdelta = -1.140881238e-8   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.914995200e-01 wkt1 = -2.940415562e-8   kt2 = -0.055045   at = 2.869166035e+05 wat = -1.246736198e-2   ute = -0.29175   ua1 = 6.8217e-10   ub1 = -1.5013e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.703840235e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.635043363e-07 wvth0 = 5.126066980e-08 pvth0 = -4.799014046e-14   k1 = 0.64774   k2 = -5.617500129e-02 lk2 = 4.181313783e-08 wk2 = 1.569135093e-08 pk2 = -2.867342818e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.824985027e-09 lua = -1.608578060e-16 wua = -1.121474495e-17 pua = -2.347394857e-22   ub = 2.914554195e-18 lub = -3.263494810e-25 wub = -5.657918221e-26 pub = 9.741688656e-31   uc = 5.912933226e-11 wuc = 5.375079648e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 3.037702044e-03 lu0 = -1.636848358e-09 wu0 = -4.804167407e-10 pu0 = 1.668986006e-15   a0 = 1.858357856e+00 la0 = 1.683195430e-07 wa0 = -4.702371158e-07 pa0 = 5.702056847e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.658669565e-01 lags = 2.613393475e-07 wags = -1.377107253e-07 pags = 1.297287768e-13   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.767954761e-03 lpdiblc2 = -7.918431740e-10 wpdiblc2 = -4.490334099e-09 ppdiblc2 = 2.584364368e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.901431008e-02 ldelta = 4.376675113e-08 wdelta = -1.560184733e-08 pdelta = 3.352079856e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.916488307e-01 lkt1 = 1.193649236e-09 wkt1 = -5.876714543e-08 pkt1 = 2.347394857e-13   kt2 = -0.055045   at = 3.018023378e+05 lat = -1.190025141e-01 wat = -2.491726966e-02 pat = 9.952954194e-8   ute = -4.502977220e-01 lute = 1.267493909e-6   ua1 = 6.682694880e-10 lua1 = 1.111262531e-16   ub1 = -1.537629899e-19 lub1 = 2.904357429e-26 wub1 = -7.336489818e-26 pub1 = 5.865083420e-31   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.407785307e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.524815609e-08 wvth0 = 5.395326185e-08 pvth0 = -5.874543012e-14   k1 = 0.64774   k2 = -4.215464154e-02 lk2 = -1.418978714e-08 wk2 = 9.740546259e-09 pk2 = -4.903534004e-15   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.840698611e-09 lua = -9.809146598e-17 wua = -1.432864504e-16 pua = 2.928077343e-22   ub = 2.803138174e-18 lub = 1.186906738e-25 wub = 2.760029889e-25 pub = -3.542973585e-31   uc = 7.363920701e-11 luc = -5.795824370e-17 wuc = -8.917843455e-18 puc = 5.709165204e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.687485181e-03 lu0 = -2.379421229e-10 wu0 = -2.259049025e-10 pu0 = 6.523639198e-16   a0 = 2.173045338e+00 la0 = -1.088668135e-06 wa0 = -4.852768404e-07 pa0 = 6.302803605e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.386443858e-01 lags = -2.936281621e-08 wags = -1.732552957e-07 pags = 2.717080090e-13   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 7.195206015e-06 lpdiblc2 = 1.023573479e-08 wpdiblc2 = 5.542977376e-12 ppdiblc2 = 7.885312286e-15   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.213994084e-02 ldelta = 7.122573161e-08 wdelta = 8.975747882e-09 pdelta = -6.465194774e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.59135   kt2 = -0.055045   at = 3.038306520e+05 lat = -1.271044123e-1   ute = -1.434315642e-01 lute = 4.174772792e-08 wute = 3.119842072e-08 pute = -1.246189717e-13   ua1 = 6.9609e-10   ub1 = -1.710349202e-19 lub1 = 9.803457293e-26 wub1 = 1.467297964e-25 pub1 = -2.926379059e-31   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos  lmin = 1.5e-06 lmax = 2e-06 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.813067111e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.336244111e-08 wvth0 = -1.173614650e-08 pvth0 = 7.226552589e-14   k1 = 0.64774   k2 = -3.363371117e-02 lk2 = -3.118393067e-08 wk2 = -8.120064724e-09 pk2 = 3.071766854e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.889882058e-09 wua = 3.528498675e-18   ub = 2.862650144e-18 wub = 9.835690056e-26   uc = 4.457871578e-11 wuc = 1.970813531e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.441714806e-03 lu0 = 2.522223145e-10 wu0 = 2.257672828e-10 pu0 = -2.484510865e-16   a0 = 2.067482699e+00 la0 = -8.781340074e-07 wa0 = -6.029682700e-07 pa0 = 8.650041477e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.529247686e-01 lags = 5.404763882e-07 wags = 2.299252068e-07 pags = -5.323951853e-13   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.782923056e-03 lpdiblc2 = 1.380594665e-08 wpdiblc2 = 1.077812241e-08 ppdiblc2 = -1.359952014e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 6.821660907e-02 ldelta = -4.061357551e-08 wdelta = -4.350031964e-08 pdelta = 4.000632133e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -0.59135   kt2 = -0.055045   at = 3.364990924e+05 lat = -1.922583498e-01 wat = -9.495773312e-02 pat = 1.893837029e-7   ute = -1.224990893e-01 wute = -3.128602158e-8   ua1 = 6.9609e-10   ub1 = -1.2188e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos  lmin = 1e-06 lmax = 1.5e-06 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.643340974e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.872631491e-08 wvth0 = -8.281899669e-08 pvth0 = 1.784917372e-13   k1 = 0.64774   k2 = -5.645174755e-02 lk2 = 2.915342883e-09 wk2 = -1.511068737e-10 pk2 = 1.880885793e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.206603053e-09 lua = 4.733078560e-16 wua = 3.155138821e-16 pua = -4.662309569e-22   ub = 2.755493369e-18 lub = 1.601350853e-25 wub = 2.039114679e-25 pub = -1.577407455e-31   uc = -5.239965021e-11 luc = 1.449244701e-16 wuc = 1.152364808e-16 puc = -1.427575595e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 4.500013503e-04 lu0 = 3.228638902e-09 wu0 = 2.186638826e-09 pu0 = -3.178777521e-15   a0 = 1.862580881e+00 la0 = -5.719287314e-07 wa0 = -2.652788887e-07 pa0 = 3.603611364e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.688342294e-01 lags = 2.178212901e-07 wags = -7.142318800e-08 pags = -8.206014406e-14   b0 = 0.0   b1 = 2.1073e-24   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {-1.699103047e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.330880713e-06 wnfactor = 4.173060348e-06 pnfactor = -6.236221385e-12   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 3.452987237e-03 lpdiblc2 = 5.981402313e-09 wpdiblc2 = -1.124546971e-08 ppdiblc2 = 1.931253593e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.891008018e-03 ldelta = 5.700900270e-08 wdelta = -2.362416664e-08 pdelta = 1.030339828e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.276895105e-01 lkt1 = -9.513423545e-08 wkt1 = -1.192971288e-08 pkt1 = 1.782776293e-14   kt2 = -9.336122080e-02 lkt2 = 5.725976036e-8   at = 2.299094310e+05 lat = -3.297075991e-02 wat = 1.583197130e-01 pat = -1.891141126e-7   ute = 5.937751710e-01 lute = -1.070400255e-06 wute = -7.278584479e-07 pute = 1.040957834e-12   ua1 = 8.047580320e-10 lua1 = -1.623935070e-16   ub1 = -3.425174720e-19 lub1 = 3.297206382e-25   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.780726907e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.437534228e-08 wvth0 = 1.051285223e-07 pvth0 = -8.403275717e-15   k1 = 0.64774   k2 = -5.238211477e-02 lk2 = -1.131499952e-09 wk2 = 1.999759504e-08 pk2 = -1.227011250e-15   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.238143166e+05 lvsat = -5.401244379e-05 wvsat = 1.863493020e-02 pvsat = -1.853057459e-8   ua = -2.705835824e-09 lua = -2.465507672e-17 wua = -1.388052570e-16 pua = -1.445600502e-23   ub = 2.955490879e-18 lub = -3.874243903e-26 wub = -7.101691666e-26 pub = 1.156480401e-31   uc = 1.177368754e-10 luc = -2.425929097e-17 wuc = -4.480754372e-17 puc = 1.639021849e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 4.002733598e-03 lu0 = -3.041980452e-10 wu0 = -1.266299825e-09 pu0 = 2.548246741e-16   a0 = 8.076930383e-01 la0 = 4.770517396e-07 wa0 = 7.871910729e-07 pa0 = -6.862149934e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 8.428720172e-01 lags = -2.535618861e-07 wags = -2.350206177e-07 pags = 8.062113999e-14   b0 = 1.567506541e-06 lb0 = -1.558728504e-12 wb0 = -1.436732679e-12 pb0 = 1.428686976e-18   b1 = 5.445233443e-08 lb1 = -5.414740135e-14 wb1 = -1.625428320e-13 pb1 = 1.616325921e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {4.667430253e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.098280545e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -2.138041016e-02 lpdiblc2 = 3.067573269e-08 wpdiblc2 = 7.611773787e-09 ppdiblc2 = 5.608929947e-16   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 5.188371922e-02 ldelta = 8.290650686e-09 wdelta = -1.973334761e-08 pdelta = 6.434367834e-15   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.790899508e-01 lkt1 = -4.402163762e-08 wkt1 = -1.714511620e-08 pkt1 = 2.301395999e-14   kt2 = -2.075418400e-02 lkt2 = -1.494067703e-8   at = 3.280447319e+05 lat = -1.305565031e-01 wat = -6.017973988e-02 pat = 2.816174338e-8   ute = -4.331209124e-01 lute = -4.925478926e-08 wute = 3.438932441e-07 pute = -2.479204861e-14   ua1 = 3.894048800e-10 lua1 = 2.506336673e-16   ub1 = 6.062986240e-19 lub1 = -6.137820877e-25 wub1 = -7.461634063e-41 pub1 = -1.094764425e-47   uc1 = -2.284941472e-11 luc1 = 1.281623960e-17   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos  lmin = 3.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 3.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-5.458335523e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.787631223e-08 wvth0 = 2.272095801e-07 pvth0 = -6.876015069e-14   k1 = 0.64774   k2 = -9.288085283e-02 lk2 = 1.889107615e-08 wk2 = 3.475633437e-08 pk2 = -8.523731978e-15   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.027510387e+05 lvsat = 1.035967218e-02 wvsat = 6.114509478e-03 pvsat = -1.234047859e-8   ua = -2.321180996e-09 lua = -2.148284235e-16 wua = -5.056044559e-16 pua = 1.668895189e-22   ub = 2.016844244e-18 lub = 4.253244576e-25 wub = 5.068723631e-25 pub = -1.700604198e-31   uc = 1.174942768e-10 luc = -2.413935022e-17 wuc = -5.975131428e-17 puc = 2.377841866e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 3.487838784e-03 lu0 = -4.963404919e-11 wu0 = -1.345330520e-09 pu0 = 2.938974495e-16   a0 = 2.037631515e+00 la0 = -1.310298433e-07 wa0 = -8.618495389e-07 pa0 = 1.290706850e-13   keta = -1.172621950e-02 lketa = -4.221090809e-10 wketa = -2.548575784e-09 pketa = 1.260015868e-15   a1 = 0.0   a2 = 0.46703705   ags = 3.300041246e-01 wags = -7.195196881e-8   b0 = -5.423438130e-06 lb0 = 1.897594541e-12 wb0 = 5.381391191e-12 pb0 = -1.942193465e-18   b1 = 5.127462474e-08 lb1 = -5.257634168e-14 wb1 = -1.530572160e-13 pb1 = 1.569429036e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {4.667430253e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.098280545e-6   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -9.666541752e-02 lpdiblc2 = 6.789664033e-08 wpdiblc2 = 4.765677346e-08 ppdiblc2 = -1.923735485e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -1.535133613e-02 ldelta = 4.153166205e-08 wdelta = 9.840399425e-08 pdelta = -5.197273398e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.776655255e-01 lkt1 = 4.714126516e-09 wkt1 = 1.455152853e-08 pkt1 = 7.343138832e-15   kt2 = -7.256047259e-02 lkt2 = 1.067235205e-08 wkt2 = 9.898600835e-08 pkt2 = -4.893868253e-14   at = 1.510890536e+05 lat = -4.306961576e-02 wat = -5.007351278e-03 pat = 8.845144503e-10   ute = -6.305393711e-01 lute = 4.834889671e-08 wute = 3.398919266e-07 pute = -2.281379724e-14   ua1 = 7.005119767e-10 lua1 = 9.682231872e-17 wua1 = 5.845858998e-16 pua1 = -2.890192689e-22   ub1 = -3.029774256e-19 lub1 = -1.642360088e-25 wub1 = -1.238000224e-24 pub1 = 6.120673106e-31   uc1 = 3.352294451e-11 luc1 = -1.505425481e-17 wuc1 = -9.089335194e-17 puc1 = 4.493767320e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.44e-6   sbref = 1.44e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.347807959e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.033336706e-8   k1 = 0.64774   k2 = -5.090782910e-02 wk2 = 1.206834424e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.714727941e-09 wua = -1.690067132e-16   ub = 2.777107609e-18 wub = 1.604568241e-25   uc = 6.996144891e-11 wuc = -5.295075195e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.894566623e-03 wu0 = -3.323400480e-10   a0 = 1.177846303e+00 wa0 = 2.921649386e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 2.878571328e-01 wags = -1.243833191e-8   b0 = 9.975197113e-08 wb0 = -9.826047966e-14   b1 = -2.427691125e-07 wb1 = 2.391392288e-13   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.532779657e-03 wpdiblc2 = -1.123525710e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.211393996e-02 wdelta = 7.812022019e-10   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.580954364e-01 wkt1 = -6.230878132e-8   kt2 = -0.055045   at = 2.648074853e+05 wat = 9.311180667e-3   ute = -2.986818441e-01 wute = 6.828199156e-9   ua1 = 6.8217e-10   ub1 = -1.5013e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.347807959e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = 3.033336706e-8   k1 = 0.64774   k2 = -5.090782910e-02 wk2 = 1.206834424e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.714727941e-09 wua = -1.690067132e-16   ub = 2.777107609e-18 wub = 1.604568241e-25   uc = 6.996144891e-11 wuc = -5.295075195e-18   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.894566623e-03 wu0 = -3.323400480e-10   a0 = 1.177846303e+00 wa0 = 2.921649386e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 2.878571328e-01 wags = -1.243833191e-8   b0 = 9.975197113e-08 wb0 = -9.826047966e-14   b1 = -2.427691125e-07 wb1 = 2.391392288e-13   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 2.532779657e-03 wpdiblc2 = -1.123525710e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.211393996e-02 wdelta = 7.812022019e-10   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.580954364e-01 wkt1 = -6.230878132e-8   kt2 = -0.055045   at = 2.648074853e+05 wat = 9.311180667e-3   ute = -2.986818441e-01 wute = 6.828199156e-9   ua1 = 6.8217e-10   ub1 = -1.5013e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.523512713e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.404654087e-07 wvth0 = 3.349754335e-08 pvth0 = -2.529569095e-14   k1 = 0.64774   k2 = -5.105819348e-02 lk2 = 1.202073004e-09 wk2 = 1.065104963e-08 pk2 = 1.133042001e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.653280831e-09 lua = -4.912327788e-16 wua = -1.803516197e-16 pua = 9.069572049e-23   ub = 2.632245133e-18 lub = 1.158088580e-24 wub = 2.215087951e-25 pub = -4.880738773e-31   uc = 6.354273773e-11 luc = 5.131374465e-17 wuc = 1.027663415e-18 puc = -5.054650154e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.753211559e-03 lu0 = 1.130048925e-09 wu0 = -2.001799574e-10 pu0 = -1.056540628e-15   a0 = 9.322933621e-01 la0 = 1.963048428e-06 wa0 = 4.419808616e-07 pa0 = -1.197688414e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 1.488204165e-01 lags = 1.111515125e-06 wags = 7.609053483e-08 pags = -7.077351723e-13   b0 = 2.337809434e-08 lb0 = 6.105633206e-13 wb0 = -2.302854508e-14 pb0 = -6.014341778e-19   b1 = -2.450250414e-07 lb1 = 1.803479742e-14 wb1 = 2.413614269e-13 pb1 = -1.776514113e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -1.294702722e-03 lpdiblc2 = 3.059842513e-08 wpdiblc2 = -4.884214698e-10 ppdiblc2 = -5.077277334e-15   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -3.869901880e-03 ldelta = 1.277812252e-07 wdelta = 6.940199893e-09 pdelta = -4.923749114e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.880771831e-01 lkt1 = 2.396860752e-07 wkt1 = -6.228538976e-08 pkt1 = -1.870014855e-16   kt2 = -0.055045   at = 2.543498940e+05 lat = 8.360216782e-02 wat = 2.182566515e-02 pat = -1.000457948e-7   ute = -4.199426246e-01 lute = 9.694071834e-07 wute = -2.990122802e-08 pute = 2.936297326e-13   ua1 = 6.682694880e-10 lua1 = 1.111262531e-16   ub1 = -2.875736061e-19 lub1 = 1.098779165e-24 wub1 = 5.844498170e-26 pub1 = -4.672325617e-31   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.941652697e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -9.195275628e-08 wvth0 = 8.036962248e-09 pvth0 = 7.640405420e-14   k1 = 0.64774   k2 = -4.036565549e-02 lk2 = -4.150820077e-08 wk2 = 7.978309123e-09 pk2 = 2.200641471e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.897261180e-09 lua = 4.833223284e-16 wua = -8.756960455e-17 pua = -2.799127610e-22   ub = 3.077949920e-18 lub = -6.222346207e-25 wub = 5.300228552e-27 pub = 3.755496210e-31   uc = 7.638915888e-11 wuc = -1.162667805e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.848898575e-03 lu0 = 7.478367087e-10 wu0 = -3.849048426e-10 pu0 = -3.186755467e-16   a0 = 1.669704516e+00 la0 = -9.824666848e-07 wa0 = 1.053802933e-08 pa0 = 5.256668347e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.880229570e-01 lags = 1.560444972e-07 wags = -1.233907585e-07 pags = 8.907290577e-14   b0 = 2.274418517e-07 lb0 = -2.045489517e-13 wb0 = -2.240411411e-13 pb0 = 2.014905358e-19   b1 = -2.396919112e-07 lb1 = -3.267857761e-15 wb1 = 2.361080377e-13 pb1 = 3.218996752e-21   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 1.212501191e-03 lpdiblc2 = 2.058364982e-08 wpdiblc2 = -1.181741272e-09 ppdiblc2 = -2.307880715e-15   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 3.276109190e-02 ldelta = -1.853761633e-08 wdelta = -1.133707573e-08 pdelta = 2.376925862e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.280716565e-01 wkt1 = -6.233220568e-8   kt2 = -0.055045   at = 3.008993547e+05 lat = -1.023349977e-01 wat = 2.887468569e-03 pat = -2.439906233e-8   ute = -1.307996642e-01 lute = -1.855454574e-07 wute = 1.875539293e-08 pute = 9.927572590e-14   ua1 = 6.9609e-10   ub1 = 9.658631218e-20 lub1 = -4.357092130e-25 wub1 = -1.168899634e-25 pub1 = 2.331253430e-31   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos  lmin = 1.5e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.402707431e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = 4.634625537e-8   k1 = 0.64774   k2 = -6.117803052e-02 wk2 = 1.901241196e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -2.654921465e-09 wua = -2.279189633e-16   ub = 2.765959035e-18 wub = 1.936022848e-25   uc = 7.638915888e-11 wuc = -1.162667805e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 3.223866840e-03 wu0 = -5.446900144e-10   a0 = 1.177091858e+00 wa0 = 2.741094467e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 4.662642812e-01 wags = -7.872925339e-8   b0 = 1.248802032e-07 wb0 = -1.230129944e-13   b1 = -2.413304279e-07 wb1 = 2.377220554e-13   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 1.153322412e-02 wpdiblc2 = -2.338921735e-9   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.346625820e-02 wdelta = 5.809239762e-10   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -5.280716565e-01 wkt1 = -6.233220568e-8   kt2 = -0.055045   at = 2.495881845e+05 wat = -9.346317198e-3   ute = -2.238328859e-01 wute = 6.853263215e-8   ua1 = 6.9609e-10   ub1 = -1.2188e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos  lmin = 1e-06 lmax = 1.5e-06 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-5.932775357e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.286533508e-07 wvth0 = 1.427012793e-07 pvth0 = -1.439929477e-13   k1 = 0.64774   k2 = -1.153577372e-01 lk2 = 8.096615360e-08 wk2 = 5.787412039e-08 pk2 = -5.807493707e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 5.213874296e+04 lvsat = 1.070308065e-01 wvsat = 7.055037601e-02 pvsat = -1.054304819e-7   ua = -1.915487792e-09 lua = -1.105009680e-15 wua = -9.562966236e-16 pua = 1.088487576e-21   ub = 1.970246112e-18 lub = 1.189113391e-24 wub = 9.774177076e-25 pub = -1.171333768e-30   uc = 1.198636970e-10 luc = -6.496834977e-17 wuc = -5.445118488e-17 puc = 6.399694301e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 4.937686227e-03 lu0 = -2.561131692e-09 wu0 = -2.233946186e-09 pu0 = 2.524424423e-15   a0 = 6.019258173e-01 la0 = 8.595281315e-07 wa0 = 9.765268607e-07 pa0 = -1.049692584e-12   keta = -1.079467086e-02 lketa = -2.667995871e-09 wketa = -1.758634901e-09 pketa = 2.628103996e-15   a1 = 0.0   a2 = 0.46703705   ags = 6.260080992e-01 lags = -2.387211616e-07 wags = -3.247517941e-07 pags = 3.676560849e-13   b0 = 3.134275134e-07 lb0 = -2.817651003e-13 wb0 = -3.087411452e-13 pb0 = 2.775521485e-19   b1 = 9.097726002e-08 lb1 = -4.966006089e-13 wb1 = -8.961696803e-14 pb1 = 4.891754365e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 4.858378491e-03 lpdiblc2 = 9.974889315e-09 wpdiblc2 = -1.262984755e-08 ppdiblc2 = 1.537875954e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -5.925143684e-02 ldelta = 1.236133235e-07 wdelta = 3.758912439e-08 pdelta = -5.530505469e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -2.582625170e-01 lkt1 = -4.032027781e-07 wkt1 = -2.773282340e-07 pkt1 = 3.212900647e-13   kt2 = -2.105544821e-01 lkt2 = 2.323933701e-07 wkt2 = 1.154409877e-07 pkt2 = -1.725150120e-13   at = 2.918183708e+05 lat = -6.310879036e-02 wat = 9.733643574e-02 pat = -1.594267060e-7   ute = -2.139097634e-01 lute = -1.482911439e-08 wute = 6.774998138e-08 pute = 1.169593302e-15   ua1 = 9.979992208e-10 lua1 = -4.511731395e-16 wua1 = -1.903518465e-16 pua1 = 2.844617994e-22   ub1 = -5.388043613e-19 lub1 = 6.230517656e-25 wub1 = 1.933520078e-25 pub1 = -2.889452404e-31   uc1 = 8.453375214e-11 luc1 = -1.412129576e-16 wuc1 = -9.308186660e-17 puc1 = 1.391015414e-22   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.019187402e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.836616461e-08 wvth0 = 3.011322573e-08 pvth0 = -3.203538728e-14   k1 = 0.64774   k2 = -2.920573114e-02 lk2 = -4.703401191e-09 wk2 = -2.832255306e-09 pk2 = 2.291482921e-15   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.863063691e+05 lvsat = -2.638548087e-02 wvsat = -4.292274108e-02 pvsat = 7.407185722e-9   ua = -3.101914627e-09 lua = 7.477316359e-17 wua = 2.513513751e-16 pua = -1.123975943e-22   ub = 3.331728366e-18 lub = -1.647445622e-25 wub = -4.416289008e-25 pub = 2.397661796e-31   uc = 6.494258832e-11 luc = -1.035479929e-17 wuc = 7.197363225e-18 puc = 2.693626773e-24   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.463957687e-03 lu0 = -1.012560321e-10 wu0 = 2.494683082e-10 pu0 = 5.491704999e-17   a0 = 1.766488568e+00 la0 = -2.985130682e-07 wa0 = -1.572685465e-07 pa0 = 7.775356940e-14   keta = -1.347769164e-02 wketa = 8.842693590e-10   a1 = 0.0   a2 = 0.46703705   ags = 7.992175134e-01 lags = -4.109606030e-07 wags = -1.920188360e-07 pags = 2.356664313e-13   b0 = 8.752903572e-08 lb0 = -5.713165414e-14 wb0 = 2.111620238e-14 pb0 = -5.045799788e-20   b1 = -5.701314862e-07 lb1 = 1.608059283e-13 wb1 = 4.527022113e-13 pb1 = -5.010675540e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = 1.300374711e-02 lpdiblc2 = 1.875134762e-09 wpdiblc2 = -2.625827157e-08 ppdiblc2 = 2.893086438e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 3.609779515e-02 ldelta = 2.879804718e-08 wdelta = -4.183454679e-09 pdelta = -1.376640207e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.582333260e-01 lkt1 = -5.471805645e-09 wkt1 = 6.081490721e-08 pkt1 = -1.495947489e-14   kt2 = 5.603687518e-02 lkt2 = -3.270507562e-08 wkt2 = -7.564287926e-08 pkt2 = 1.749878530e-14   at = 4.406018237e+05 lat = -2.110590560e-01 wat = -1.710538781e-01 pat = 1.074606221e-7   ute = -6.499298767e-02 lute = -1.629119561e-07 wute = -1.873043193e-08 pute = 8.716571630e-14   ua1 = -7.440364279e-12 lua1 = 5.486359839e-16 wua1 = 3.909116142e-16 pua1 = -2.935465859e-22   ub1 = 1.221374061e-18 lub1 = -1.127269657e-24 wub1 = -6.058788287e-25 pub1 = 5.058099033e-31   uc1 = -8.568713394e-11 luc1 = 2.805469152e-17 wuc1 = 6.189816964e-17 puc1 = -1.501060659e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos  lmin = 3.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 1.0e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.782289999e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -7.222604304e-08 wvth0 = -1.348985490e-07 pvth0 = 4.954643417e-14   k1 = 0.64774   k2 = -4.695523411e-02 lk2 = 4.071953082e-09 wk2 = -1.048260450e-08 pk2 = 6.073815561e-15   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.729186447e+05 lvsat = -1.976658997e-02 wvsat = -6.300395056e-02 pvsat = 1.733533569e-8   ua = -3.076683126e-09 lua = 6.229870963e-17 wua = 2.386014056e-16 pua = -1.060940094e-22   ub = 2.612994519e-18 lub = 1.905974519e-25 wub = -8.036427329e-26 pub = 6.115694775e-32   uc = 1.607392219e-11 luc = 1.380586924e-17 wuc = 4.015260322e-17 puc = -1.359944388e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 9.335311068e-04 lu0 = 6.553868693e-10 wu0 = 1.170785149e-09 pu0 = -4.005819962e-16   a0 = 1.1627   keta = -1.727227166e-02 lketa = 1.876040360e-09 wketa = 2.914551807e-09 pketa = -1.003771642e-15   a1 = 0.0   a2 = 0.46703705   ags = -7.446080985e-01 lags = 3.523067795e-07 wags = 9.865926523e-07 pags = -3.470390885e-13   b0 = 7.894683512e-07 lb0 = -4.041704517e-13 wb0 = -7.386199123e-13 pb0 = 3.251555372e-19   b1 = -1.841702328e-06 lb1 = 7.894705525e-13 wb1 = 1.711615945e-12 pb1 = -6.725137054e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = 0.030097   pdiblc1 = 0.0   pdiblc2 = -2.703778191e-03 lpdiblc2 = 9.640935270e-09 wpdiblc2 = -4.489995143e-08 ppdiblc2 = 3.814731091e-14   pdiblcb = -0.025   drout = 0.43496   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.509909476e-01 ldelta = -2.800512739e-08 wdelta = -6.545113965e-08 pdelta = 1.652434138e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -7.924373247e-01 lkt1 = 6.087865133e-08 wkt1 = 1.276072598e-07 pkt1 = -4.798161401e-14   kt2 = 1.626020472e-01 lkt2 = -8.539089664e-08 wkt2 = -1.326603614e-07 pkt2 = 4.568822846e-14   at = -4.433949910e+04 lat = 2.869593405e-02 wat = 1.874991537e-01 pat = -6.980799686e-8   ute = -8.127409949e-01 lute = 2.067746586e-07 wute = 5.193692717e-07 pute = -1.788707772e-13   ua1 = 1.972651465e-09 lua1 = -4.303214166e-16 wua1 = -6.685325589e-16 pua1 = 2.302426133e-22   ub1 = -2.955731024e-18 lub1 = 9.378910967e-25 wub1 = 1.375089403e-24 pub1 = -4.735807904e-31   uc1 = -1.642735167e-10 luc1 = 6.690779914e-17 wuc1 = 1.039456565e-16 puc1 = -3.579888411e-23   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.44e-6   sbref = 1.44e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos  lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.478440006e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = -1.618199141e-8   k1 = 0.64774   k2 = -2.013907286e-02 wk2 = -4.394417249e-9   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.354638400e-09 wua = 1.733760978e-16   ub = 3.679898369e-18 wub = -3.225795667e-25   uc = 5.987805477e-11 wuc = 1.000246718e-19   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.061043755e-03 wu0 = 1.136346955e-10   a0 = 2.042018468e+00 wa0 = -1.702086499e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 6.141664240e-01 wags = -1.870294655e-7   b0 = 6.018892086e-08 wb0 = -7.709234874e-14   b1 = 1.270027772e-07 wb1 = 4.129351869e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -4.524491454e-01 wpclm = 2.581853500e-7   pdiblc1 = 0.0   pdiblc2 = 1.367614996e-03 wpdiblc2 = -5.001066884e-10   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.031492148e-02 wdelta = 1.743763446e-9   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -8.614952308e-01 wkt1 = 1.000246718e-7   kt2 = -0.055045   at = 2.574397569e+05 wat = 1.325326902e-2   ute = -6.244466554e-01 wute = 1.811280099e-7   ua1 = 6.8217e-10   ub1 = -7.061596185e-20 wub1 = -4.254382709e-26   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos  lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.243608117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.695322724e-07 wvth0 = -2.874662467e-08 pvth0 = 2.512223033e-13   k1 = 0.64774   k2 = -1.514593992e-02 lk2 = -9.983469732e-08 wk2 = -7.065983044e-09 pk2 = 5.341635513e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.354638400e-09 wua = 1.733760978e-16   ub = 3.679898369e-18 wub = -3.225795667e-25   uc = 5.987805477e-11 wuc = 1.000246718e-19   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.136018588e-03 lu0 = -1.499076810e-09 wu0 = 7.351956082e-11 pu0 = 8.020780492e-16   a0 = 1.691430168e+00 la0 = 7.009802693e-06 wa0 = 1.737291849e-08 pa0 = -3.750580911e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 6.141664240e-01 wags = -1.870294655e-7   b0 = 2.194793063e-07 lb0 = -3.184915682e-12 wb0 = -1.623203509e-13 pb0 = 1.704082766e-18   b1 = 1.229343754e-07 lb1 = 8.134525327e-14 wb1 = 4.347030894e-14 pb1 = -4.352361507e-20   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -4.524491454e-01 wpclm = 2.581853500e-7   pdiblc1 = 0.0   pdiblc2 = 3.630289878e-03 lpdiblc2 = -4.524082665e-08 wpdiblc2 = -1.710746358e-09 ppdiblc2 = 2.420601382e-14   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.189948808e-02 ldelta = -2.316264584e-07 wdelta = -4.454535745e-09 pdelta = 1.239312733e-13   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -8.614952308e-01 wkt1 = 1.000246718e-7   kt2 = -0.055045   at = 2.233565131e+05 lat = 6.814740096e-01 wat = 3.148944044e-02 pat = -3.646213059e-7   ute = -6.244466554e-01 wute = 1.811280099e-7   ua1 = 6.8217e-10   ub1 = -1.764370963e-20 lub1 = -1.059148400e-24 wub1 = -7.088652469e-26 pub1 = 5.666952330e-31   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos  lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-4.492072512e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.285401037e-07 wvth0 = 3.181534166e-08 pvth0 = -2.329342803e-13   k1 = 0.64774   k2 = -4.463150842e-02 lk2 = 1.358847315e-07 wk2 = 7.212464642e-09 pk2 = -6.073126705e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.406803156e-09 lua = 4.170259269e-16 wua = 2.228189933e-16 pua = -3.952662835e-22   ub = 4.024686478e-18 lub = -2.756374060e-24 wub = -5.235141620e-25 pub = 1.606351529e-30   uc = 1.008054692e-10 luc = -3.271901221e-16 wuc = -1.890968655e-17 puc = 1.519712354e-22   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.686015463e-03 lu0 = -5.895971827e-09 wu0 = -1.642268209e-10 pu0 = 2.702717723e-15   a0 = 2.920394094e+00 la0 = -2.815026516e-06 wa0 = -6.217484589e-07 pa0 = 1.358811028e-12   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 7.229168068e-01 lags = -8.693940601e-07 wags = -2.310785906e-07 pags = 3.521463253e-13   b0 = -1.298512293e-07 lb0 = -3.922276485e-13 wb0 = 5.895649806e-14 pb0 = -6.489287536e-20   b1 = 2.069423730e-07 lb1 = -5.902482824e-13 wb1 = -4.628341615e-16 pb1 = 3.076955042e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -4.524491454e-01 wpclm = 2.581853500e-7   pdiblc1 = 0.0   pdiblc2 = 1.563549316e-03 lpdiblc2 = -2.871847591e-08 wpdiblc2 = -2.017723507e-09 ppdiblc2 = 2.666011193e-14   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -4.113715150e-03 ldelta = -2.366650655e-08 wdelta = 7.070651696e-09 pdelta = 3.179431485e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -9.847750125e-01 lkt1 = 9.855478870e-07 wkt1 = 1.499669905e-07 pkt1 = -3.992588722e-13   kt2 = -0.055045   at = 3.478857935e+05 lat = -3.140628697e-01 wat = -2.822053080e-02 pat = 1.127240882e-7   ute = -1.152407130e+00 lute = 4.220727217e-06 wute = 3.620024406e-07 pute = -1.445982549e-12   ua1 = 6.682694880e-10 lua1 = 1.111262531e-16   ub1 = -1.783404500e-19 lub1 = 2.255256215e-25   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos  lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.566101092e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.586700798e-07 wvth0 = -1.205685125e-08 pvth0 = -5.769119301e-14   k1 = 0.64774   k2 = -1.521082292e-02 lk2 = 1.836674536e-08 wk2 = -5.480733731e-09 pk2 = -1.002955547e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.261358213e-09 lua = -1.639393526e-16 wua = 1.072397848e-16 pua = 6.640330687e-23   ub = 3.252542285e-18 lub = 3.278787051e-25 wub = -8.811506757e-26 pub = -1.328066137e-31   uc = 1.889326160e-11 wuc = 1.913638680e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.207947312e-03 lu0 = 8.023598006e-12 wu0 = 4.930828488e-10 pu0 = 7.715997855e-17   a0 = 2.005615615e+00 la0 = 8.389646433e-07 wa0 = -1.691905321e-07 pa0 = -4.488863545e-13   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 3.434268171e-01 lags = 6.464407545e-07 wags = -9.952968307e-08 pags = -1.733126309e-13   b0 = -3.687375558e-07 lb0 = 5.619798943e-13 wb0 = 9.494345851e-14 pb0 = -2.086391902e-19   b1 = -6.948688381e-09 lb1 = 2.641181731e-13 wb1 = 1.115792419e-13 pb1 = -1.398453643e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -4.524491454e-01 wpclm = 2.581853500e-7   pdiblc1 = 0.0   pdiblc2 = -1.691889235e-02 lpdiblc2 = 4.510778909e-08 wpdiblc2 = 8.519424580e-09 ppdiblc2 = -1.542947238e-14   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = -4.848766842e-02 ldelta = 1.535808124e-07 wdelta = 3.213491098e-08 pdelta = -6.832236244e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -6.927731921e-01 lkt1 = -1.808241842e-07 wkt1 = 2.579102155e-08 pkt1 = 9.674961811e-14   kt2 = -0.055045   at = 3.062960080e+05 lat = -1.479366304e-1   ute = -1.433581237e-01 lute = 1.901818668e-07 wute = 2.547477154e-08 pute = -1.017564275e-13   ua1 = 6.9609e-10   ub1 = -1.2188e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos  lmin = 1.5e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-2.770523074e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = -4.098344221e-8   k1 = 0.64774   k2 = -6.001664603e-03 wk2 = -1.050959227e-8   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 123760.0   ua = -3.343558049e-09 wua = 1.405346639e-16   ub = 3.416941957e-18 wub = -1.547048258e-25   uc = 1.889326160e-11 wuc = 1.913638680e-17   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 1.211970375e-03 wu0 = 5.317711653e-10   a0 = 2.426275785e+00 wa0 = -3.942639148e-7   keta = -0.01258   a1 = 0.0   a2 = 0.46703705   ags = 6.675547526e-01 wags = -1.864293175e-7   b0 = -8.695862769e-08 wb0 = -9.669051610e-15   b1 = 1.254812018e-07 wb1 = 4.146022647e-14   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -4.524491454e-01 wpclm = 2.581853500e-7   pdiblc1 = 0.0   pdiblc2 = 5.698330418e-03 wpdiblc2 = 7.830264727e-10   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 2.851835465e-02 wdelta = -2.122190121e-9   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -7.834391489e-01 wkt1 = 7.430166039e-8   kt2 = -0.055045   at = 232120.0   ute = -4.800018806e-02 wute = -2.554630119e-8   ua1 = 6.9609e-10   ub1 = -1.2188e-19   uc1 = -9.961e-12   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 3.0e-6   sbref = 3.0e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos  lmin = 1e-06 lmax = 1.5e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-2.069790807e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.047174300e-07 wvth0 = -6.398693646e-08 pvth0 = 3.437642181e-14   k1 = 0.64774   k2 = 1.968102556e-02 lk2 = -3.838021218e-08 wk2 = -1.437809953e-08 pk2 = 5.781097254e-15   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 3.716797359e+05 lvsat = -3.704912534e-01 wvsat = -1.004193932e-01 pvsat = 1.500667412e-7   ua = -4.494026749e-09 lua = 1.719260425e-15 wua = 4.233454880e-16 pua = -4.226324955e-22   ub = 5.192268265e-18 lub = -2.653047635e-24 wub = -7.465188011e-25 pub = 8.844068047e-31   uc = -7.809398269e-11 luc = 1.449377379e-16 wuc = 5.146567573e-17 puc = -4.831288937e-23   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.384305083e-04 lu0 = 1.454857977e-09 wu0 = 2.803811874e-10 pu0 = 3.756771829e-16   a0 = 4.443521928e+00 la0 = -3.014572636e-06 wa0 = -1.078911455e-06 pa0 = 1.023137284e-12   keta = -1.875998549e-02 lketa = 9.235370321e-09 wketa = 2.503190764e-09 pketa = -3.740768278e-15   a1 = 0.0   a2 = 0.46703705   ags = -9.074681559e-01 lags = 2.353714235e-06 wags = 4.957316092e-07 pags = -1.019421289e-12   b0 = -1.221855074e-06 lb0 = 1.695989250e-12 wb0 = 5.127087328e-13 pb0 = -7.806413610e-19   b1 = 2.928947411e-07 lb1 = -2.501827931e-13 wb1 = -1.976525125e-13 pb1 = 3.573300771e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -4.524491454e-01 wpclm = 2.581853500e-7   pdiblc1 = 0.0   pdiblc2 = -4.490180179e-02 lpdiblc2 = 7.561683757e-08 wpdiblc2 = 1.399423738e-08 ppdiblc2 = -1.974283358e-14   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.936825423e-02 ldelta = 1.367391006e-08 wdelta = -4.476184084e-09 pdelta = 3.517808579e-15   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -1.172057365e+00 lkt1 = 5.807510617e-07 wkt1 = 2.115958717e-07 pkt1 = -2.051724694e-13   kt2 = 5.203707200e-03 lkt2 = -9.003566804e-8   at = 9.767182471e+05 lat = -1.112727620e+00 wat = -2.691178733e-01 pat = 4.021697498e-7   ute = -1.800541895e-01 lute = 1.973414998e-07 wute = 4.963562433e-08 pute = -1.123518695e-13   ua1 = 3.733623339e-10 lua1 = 4.822842242e-16 wua1 = 1.438588705e-16 pua1 = -2.149826961e-22   ub1 = -4.568487561e-19 lub1 = 5.005773090e-25 wub1 = 1.495018251e-25 pub1 = -2.234155274e-31   uc1 = -8.943543680e-11 luc1 = 1.187665984e-16 wuc1 = -6.162975822e-33 puc1 = 1.175494351e-38   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 2.74e-6   sbref = 2.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos  lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-1.629749793e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = -1.484751085e-07 wvth0 = -9.773315568e-08 pvth0 = 6.793366220e-14   k1 = 0.64774   k2 = 1.819576475e-02 lk2 = -3.690326883e-08 wk2 = -2.819433088e-08 pk2 = 1.951995770e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = 1.353921311e+05 lvsat = -1.355268591e-01 wvsat = -1.568117988e-02 pvsat = 6.580306187e-8   ua = -2.759653720e-09 lua = -5.400115163e-18 wua = 6.822536163e-17 pua = -6.950104183e-23   ub = 2.124083669e-18 lub = 3.979551280e-25 wub = 2.045189795e-25 pub = -6.130516426e-32   uc = 8.818359686e-11 luc = -2.040868724e-17 wuc = -5.237691916e-18 puc = 8.072939411e-24   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 5.449906252e-04 lu0 = 1.150014597e-09 wu0 = 1.276207797e-09 pu0 = -6.145727974e-16   a0 = 3.281140972e+00 la0 = -1.858701013e-06 wa0 = -9.676802856e-07 pa0 = 9.125290091e-13   keta = -9.472605846e-03 wketa = -1.258643787e-9   a1 = 0.0   a2 = 0.46703705   ags = 1.337411384e+00 lags = 1.214060196e-07 wags = -4.799783903e-07 pags = -4.917526545e-14   b0 = 1.107522025e-06 lb0 = -6.203433373e-13 wb0 = -5.246290063e-13 pb0 = 2.508872868e-19   b1 = -9.415855486e-07 lb1 = 9.773844070e-13 wb1 = 6.514479645e-13 pb1 = -4.870154372e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -8.285602172e-01 lpclm = 3.740048498e-07 wpclm = 4.594228267e-07 ppclm = -2.001105469e-13   pdiblc1 = 0.0   pdiblc2 = -1.252641263e-01 lpdiblc2 = 1.555291331e-07 wpdiblc2 = 4.772167757e-08 ppdiblc2 = -5.328140011e-14   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 9.424127375e-02 ldelta = -6.077982055e-08 wdelta = -3.529300662e-08 pdelta = 3.416205691e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -4.597726427e-01 lkt1 = -1.275448658e-07 wkt1 = -4.537108445e-08 pkt1 = 5.035547182e-14   kt2 = -0.085339   at = -3.012027963e+05 lat = 1.580370651e-01 wat = 2.258472002e-01 pat = -9.002351928e-8   ute = 1.354712275e-01 lute = -1.164169749e-07 wute = -1.259884093e-07 pute = 6.228866957e-14   ua1 = 9.029117574e-10 lua1 = -4.429972254e-17 wua1 = -9.617046783e-17 pua1 = 2.370247795e-23   ub1 = 8.905531727e-19 lub1 = -8.392791689e-25 wub1 = -4.288737743e-25 pub1 = 3.517211686e-31   uc1 = 3.0e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.74e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos  lmin = 3.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 4.23e-9   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = 2.8e-9   ll = 0.0   lw = 0.0   lwl = 0.0   wint = 7.476e-9   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = -7.916e-9   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.69   rnoib = 0.34   tnoia = 25000000.0   tnoib = 0.0   epsrox = 3.9   toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7000000000000000e+17   nsd = 1.0e+20   rshg = 0.1   rsh = 1.0   vth0 = {-3.120368596e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -7.477891485e-08 wvth0 = -6.330492130e-08 pvth0 = 5.091234313e-14   k1 = 0.64774   k2 = -3.584916732e-02 lk2 = -1.018345441e-08 wk2 = -1.642488332e-08 pk2 = 1.370114283e-14   k3 = 3.39   dvt0 = 2.4422   dvt1 = 0.16136   dvt2 = 0.026237   dvt0w = 0.5   dvt1w = 1928100.0   dvt2w = -0.032   w0 = 1.0e-8   k3b = 1.0   phin = 0.0   lpe0 = 0.0   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = -4.914187452e+05 lvsat = 1.743684381e-01 wvsat = 2.924484413e-01 pvsat = -8.653622282e-8   ua = -2.073443004e-09 lua = -3.446626931e-16 wua = -2.981802150e-16 pua = 1.116498753e-22   ub = 1.320790852e-18 lub = 7.951030964e-25 wub = 6.110267143e-25 pub = -2.622825884e-31   uc = 7.979688230e-11 luc = -1.626229556e-17 wuc = 6.057760859e-18 puc = 2.488467559e-24   rdsw = 484.7   prwb = 0.1   prwg = 0.052   wr = 1.0   u0 = 2.842284075e-03 lu0 = 1.423271530e-11 wu0 = 1.495106913e-10 pu0 = -5.753374844e-17   a0 = -4.783675508e-01 wa0 = 8.780499109e-7   keta = -9.472605846e-03 wketa = -1.258643787e-9   a1 = 0.0   a2 = 0.46703705   ags = 4.049647402e+00 lags = -1.219523467e-06 wags = -1.578564165e-06 pags = 4.939655414e-13   b0 = -4.852296558e-07 lb0 = 1.671130935e-13 wb0 = -5.659529299e-14 pb0 = 1.949141890e-20   b1 = 3.412430078e-06 lb1 = -1.175240919e-12 wb1 = -1.099597091e-12 pb1 = 3.787012380e-19   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = 0.0   cit = -6.393105e-11   cdsc = 2.8125e-7   cdscb = 1.0e-4   cdscd = 1.0e-10   eta0 = 0.2   etab = -0.00025   dsub = 1.0   voffl = 0.0   minv = 0.0   pclm = -7.207791588e-02 wpclm = 5.466848439e-8   pdiblc1 = 0.0   pdiblc2 = -7.566071834e-02 lpdiblc2 = 1.310052082e-07 wpdiblc2 = -5.864486519e-09 ppdiblc2 = -2.678840058e-14   pdiblcb = -0.025   drout = 4.620670585e-01 wdrout = -1.450357742e-8   pscbe1 = 800000000.0   pscbe2 = 8.6797e-9   pvag = 0.0   delta = 1.275507657e-01 ldelta = -7.724803336e-08 wdelta = -5.290951719e-08 pdelta = 4.287165974e-14   alpha0 = 5.0449517e-13   alpha1 = -4.0583656e-18   beta0 = 6.2016506   fprout = 0.0   pdits = 0.0   pditsl = 0.0   pditsd = 0.0   agidl = 0.0   bgidl = 2300000000.0   cgidl = 0.5   egidl = 0.8   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 4.23e-9   kt1 = -9.018719761e-01 lkt1 = 9.102904455e-08 wkt1 = 1.861600511e-07 pkt1 = -6.411352160e-14   kt2 = -0.085339   at = 3.651974523e+04 lat = -8.932959457e-03 wat = 1.442355768e-01 pat = -4.967473264e-8   ute = 1.579556000e-01 lute = -1.275332486e-7   ua1 = 1.020267349e-09 lua1 = -1.023203270e-16 wua1 = -1.589613423e-16 pua1 = 5.474628630e-23   ub1 = -2.126180082e-18 lub1 = 6.521937523e-25 wub1 = 9.312398306e-25 pub1 = -3.207189977e-31   uc1 = 3.0e-11   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 3.0e+41   noib = 0.0   noic = 0.0   em = 41000000.0   af = 1.0   ef = 0.88   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.3632   jss = 2.1483e-5   jsws = 1.4472e-10   xtis = 5.2   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.001671   tpbsw = 0.001246   tpbswg = 0.0   tcj = 0.0012407   tcjsw = 0.00037357   tcjswg = 2.0e-12   cgdo = 2.0e-11   cgso = 2.0e-11   cgbo = 1.0e-13   capmod = 2.0   xpart = 0.0   cgsl = 0.0   cgdl = 0.0   cf = 0.0   clc = 7.0e-8   cle = 0.492   dlc = -1.2e-8   dwc = 0.0   vfbcv = -1.0   acde = 0.44   moin = 8.7   noff = 2.6123   voffcv = 0.112   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = 0.0007653568198   mjs = 0.3362   pbs = 0.6587   cjsws = 9.1602368e-11   mjsws = 0.2659   pbsws = 0.7418   cjswgs = 2.39155046e-10   mjswgs = 0.9274   pbswgs = 1.4338   saref = 1.44e-6   sbref = 1.44e-6   wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}   lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}   wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__pfet_01v8_lvt





















