** Translated using xdm 2.6.0 on Nov_14_2022_16_05_13_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 2
.PARAM 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__TOXE_MULT=1.042 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__RBPB_MULT=1.2 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__OVERLAP_MULT=0.99758 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__AJUNCTION_MULT=1.1193 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__PJUNCTION_MULT=1.1801 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__LINT_DIFF=-1.21275e-8 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__WINT_DIFF=2.252e-8 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__RSHG_DIFF=7.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__DLC_DIFF=-1.21275e-8 SKY130_FD_PR__RF_NFET_G5V0D10V5_B__DWC_DIFF=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_B__XGW_DIFF=4.504e-8 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VTH0_DIFF_0=0.037892 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__NFACTOR_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VSAT_DIFF_0=-7490.2 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__K2_DIFF_0=0.0061192 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__U0_DIFF_0=-0.0068374 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UB_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VTH0_DIFF_1=0.042869 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__UA_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__VSAT_DIFF_1=-5260.5 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__A0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__RDSW_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__AGS_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__K2_DIFF_1=0.0082977 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__PCLM_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__U0_DIFF_1=-0.0034898 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM02__B1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VSAT_DIFF_0=-7602.3 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VTH0_DIFF_0=0.028278 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__K2_DIFF_0=0.0058947 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__U0_DIFF_0=-0.0070921 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VSAT_DIFF_1=-7404.4 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VTH0_DIFF_1=0.035525 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__K2_DIFF_1=0.0078725 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__U0_DIFF_1=-0.0038822 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__NFACTOR_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VSAT_DIFF_2=-8487.7 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VTH0_DIFF_2=0.039934 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__A0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__K2_DIFF_2=0.0052827 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__U0_DIFF_2=-0.0061567 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__AGS_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM04__UA_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__K2_DIFF_0=0.0053572 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__U0_DIFF_0=-0.0056999 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VTH0_DIFF_0=0.037862 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VSAT_DIFF_0=86.018 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_0=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_0=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__K2_DIFF_1=0.001022 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__U0_DIFF_1=-0.0060669 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_1=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VTH0_DIFF_1=0.032656 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VSAT_DIFF_1=-8977.1 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_1=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__A0_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B0_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UA_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__RDSW_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__K2_DIFF_2=0.0043107 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__KT1_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__U0_DIFF_2=-0.011734 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__B1_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VOFF_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__NFACTOR_DIFF_2=0.0 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__UB_DIFF_2=0.0 SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VTH0_DIFF_2=0.025004 
+ SKY130_FD_PR__RF_NFET_G5V0D10V5_BM10__VSAT_DIFF_2=-884.49
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
*





* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 002, W = 7.09, L = 0.5
* --------------------------------------------
*















* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 000, W = 3.01, L = 0.5
* ---------------------------------------------
*















* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 001, W = 5.05, L = 0.5
* ---------------------------------------------
*















* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 002, W = 7.09, L = 0.5
* ---------------------------------------------
.INCLUDE sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice















