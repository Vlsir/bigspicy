** Translated using xdm 2.6.0 on Nov_14_2022_16_05_17_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TOXE_MULT=0.94 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RSHP_MULT=1.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__OVERLAP_MULT=0.70 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AJUNCTION_MULT=9.3222e-1 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PJUNCTION_MULT=9.4436e-1 SKY130_FD_PR__ESD_PFET_G5V0D10V5__LINT_DIFF=1.7325e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__WINT_DIFF=-3.2175e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__DLC_DIFF=1.7325e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__DWC_DIFF=-3.2175e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_0=-0.0038637 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_0=0.0001511 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_0=-39322.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_0=0.059104 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_0=-0.10802 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_0=2.5385e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_0=-3.7667e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_0=0.020009 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_1=0.010686 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_1=-0.0040259 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_1=0.00027138 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_1=-36371.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_1=0.06664 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_1=2.9833e-13 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_1=-0.027795 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_1=-3.4315e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_2=0.016012 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_2=-0.0035475 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_2=-2.9036e-5 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_2=0.068406 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_2=6.8019e-12 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_2=-35489.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_2=-0.067543 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_2=-3.2017e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_3=0.018257 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_3=-0.0039581 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_3=0.00037927 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_3=0.062703 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_3=7.5609e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_3=-41289.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_3=-0.086391 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_3=-3.2769e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_4=0.016385 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_4=-0.0035685 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_4=-9.8839e-5 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_4=0.059795 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_4=-3.5551e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_4=-32637.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_4=-0.066648 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_4=-3.8565e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_5=0.019428 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_5=-0.0042313 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_5=0.00026379 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_5=0.061609 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_5=3.0966e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_5=-31131.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_5=-0.1004 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_5=-2.4624e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_6=-3.0234e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_6=0.018078 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_6=-0.0038572 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_6=7.053e-5 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_6=0.063062 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_6=2.686e-12 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_6=-32971.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_6=-0.084269 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_7=-3.572e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_7=0.021219 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_7=-0.0040301 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_7=0.00017124 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_7=0.063527 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_7=-8.4538e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_7=-29165.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_7=-0.11422 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_7=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
*




* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
.INCLUDE sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice























