** Translated using xdm 2.6.0 on Nov_14_2022_16_05_25_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NFET_03V3_NVT__TOXE_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_03V3_NVT__VTH0_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_03V3_NVT__VOFF_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_SLOPE_SPECTRE=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_03v3_nvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_03v3_nvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_03v3_nvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_03v3_nvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.SUBCKT sky130_fd_pr__nfet_03v3_nvt d g s b
.PARAM L=1 W=1 NF=1.0 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 SA=0 SB=0 SD=0 MULT=1

* msky130_fd_pr__nfet_03v3_nvt d g s b sky130_fd_pr__nfet_03v3_nvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}; HSpice Parser Retained (as a comment). Continuing.
* .model sky130_fd_pr__nfet_03v3_nvt__model.0 nmos  lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.995e-06 wmax = 1.0005e-5   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {-0.0007337+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.27   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_0}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {116050+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0}   ua = {5.1975e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_0}   ub = {5.727e-020+sky130_fd_pr__nfet_03v3_nvt__ub_diff_0}   uc = 1.3541e-10   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.091551+sky130_fd_pr__nfet_03v3_nvt__u0_diff_0}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_0}   keta = {0.0070658+sky130_fd_pr__nfet_03v3_nvt__keta_diff_0}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_0}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_0}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_0}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.0354+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0.017338+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0}   etab = 0.0   dsub = 0.59286   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 6.234e-7   alpha1 = 0.0   beta0 = 21.814   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.33884+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0}   kt2 = 0.0   at = 40500.0   ute = -1.716   ua1 = 1.0e-9   ub1 = -1.18e-17   uc1 = -3.696e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.745e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.
* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.1 nmos  lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {-0.0007337+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.27   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_1}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.018557   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {125130+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1}   ua = {4.848e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_1}   ub = {5.727e-020+sky130_fd_pr__nfet_03v3_nvt__ub_diff_1}   uc = 1.3541e-10   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.087889+sky130_fd_pr__nfet_03v3_nvt__u0_diff_1}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_1}   keta = {0.019064+sky130_fd_pr__nfet_03v3_nvt__keta_diff_1}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_1}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_1}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_1}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_1+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.0354+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0.0017338+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1}   etab = 1.0e-10   dsub = 0.59286   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 4.8972e-7   alpha1 = 0.03   beta0 = 20.82   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.33884+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1}   kt2 = -0.02   at = 40500.0   ute = -1.716   ua1 = 1.0e-9   ub1 = -1.2744e-17   uc1 = -2.5133e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.745e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.2 nmos  lmin = 5.95e-07 lmax = 6.05e-07 wmin = 9.95e-07 wmax = 1.005e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {0.068092+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.33502   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_2}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {118050+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2}   ua = {4.145e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_2}   ub = {3.7798e-019+sky130_fd_pr__nfet_03v3_nvt__ub_diff_2}   uc = 1.3541e-10   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.083529+sky130_fd_pr__nfet_03v3_nvt__u0_diff_2}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_2}   keta = {-0.016684+sky130_fd_pr__nfet_03v3_nvt__keta_diff_2}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_2}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_2}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_2}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_2+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.77345+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2}   etab = 0.0   dsub = 0.071143   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 8.3952e-7   alpha1 = 0.33   beta0 = 23.0   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.29818+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2}   kt2 = -0.02   at = 37260.0   ute = -1.613   ua1 = 1.0e-9   ub1 = -8.411e-18   uc1 = -2.5133e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.95e-6   sbref = 1.94e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.3 nmos  lmin = 4.95e-07 lmax = 5.05e-07 wmin = 3.995e-06 wmax = 4.005e-6   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {-0.0007337+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.27   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_3}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {118050+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3}   ua = {5.05e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_3}   ub = {5.727e-020+sky130_fd_pr__nfet_03v3_nvt__ub_diff_3}   uc = 1.3541e-10   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.087889+sky130_fd_pr__nfet_03v3_nvt__u0_diff_3}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_3}   keta = {0.0070658+sky130_fd_pr__nfet_03v3_nvt__keta_diff_3}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_3}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_3}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_3}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_3+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.0354+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0.017338+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3}   etab = 0.0   dsub = 0.59286   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 7.6956e-7   alpha1 = 0.0   beta0 = 22.396   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.33884+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3}   kt2 = -0.02   at = 40500.0   ute = -1.716   ua1 = 1.0e-9   ub1 = -1.2744e-17   uc1 = -2.5133e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.745e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.4 nmos  lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {-0.022934+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.30326   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_4}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {133130+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4}   ua = {4.1034e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_4}   ub = {4.971e-020+sky130_fd_pr__nfet_03v3_nvt__ub_diff_4}   uc = 2.1124e-11   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.084373+sky130_fd_pr__nfet_03v3_nvt__u0_diff_4}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_4}   keta = {0.030502+sky130_fd_pr__nfet_03v3_nvt__keta_diff_4}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_4}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_4}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_4}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_4+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.0354+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0.00020806+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4}   etab = 1.0e-10   dsub = 0.59286   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 5.4233e-7   alpha1 = 0.0   beta0 = 21.174   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.35239+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4}   kt2 = -0.02   at = 40500.0   ute = -1.5444   ua1 = 1.0e-9   ub1 = -9.4306e-18   uc1 = -1.2064e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.745e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.5 nmos  lmin = 5.95e-07 lmax = 6.05e-07 wmin = 4.15e-07 wmax = 4.25e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {0.007535+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.33965   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_5}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {127800+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5}   ua = {3.7751e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_5}   ub = {4.4739e-020+sky130_fd_pr__nfet_03v3_nvt__ub_diff_5}   uc = 6.2248e-11   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.079311+sky130_fd_pr__nfet_03v3_nvt__u0_diff_5}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_5}   keta = {0.0018301+sky130_fd_pr__nfet_03v3_nvt__keta_diff_5}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_5}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_5}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_5}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_5+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.0354+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0.00020806+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5}   etab = 1.0e-10   dsub = 0.59286   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 5.3596e-7   alpha1 = 0.0   beta0 = 21.074   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.33884+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5}   kt2 = -0.02   at = 40500.0   ute = -1.5444   ua1 = 1.0e-9   ub1 = -8.6659e-18   uc1 = -2.5133e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.95e-6   sbref = 1.94e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.6 nmos  lmin = 7.95e-07 lmax = 8.05e-07 wmin = 4.15e-07 wmax = 4.25e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {0.071092+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.40202   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_6}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {117770+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6}   ua = {2.9844e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_6}   ub = {3.7798e-019+sky130_fd_pr__nfet_03v3_nvt__ub_diff_6}   uc = 7.3121e-11   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.073506+sky130_fd_pr__nfet_03v3_nvt__u0_diff_6}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_6}   keta = {0+sky130_fd_pr__nfet_03v3_nvt__keta_diff_6}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_6}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_6}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_6}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_6+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.77345+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6}   etab = 0.0   dsub = 0.071143   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 8.5632e-7   alpha1 = 0.09   beta0 = 21.989   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.30496+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6}   kt2 = -0.02   at = 28350.0   ute = -1.613   ua1 = 1.0e-9   ub1 = -6.8818e-18   uc1 = -1.3069e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 2.34e-6   sbref = 2.34e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.7 nmos  lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.95e-07 wmax = 7.05e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {-0.011467+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.2808   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_7}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {128010+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7}   ua = {4.4602e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_7}   ub = {8.0178e-020+sky130_fd_pr__nfet_03v3_nvt__ub_diff_7}   uc = 7.0413e-11   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.084373+sky130_fd_pr__nfet_03v3_nvt__u0_diff_7}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_7}   keta = {0.019064+sky130_fd_pr__nfet_03v3_nvt__keta_diff_7}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_7}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_7}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_7}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_7+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {2.0354+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0.00020806+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7}   etab = 1.0e-10   dsub = 0.59286   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 3.9877e-7   alpha1 = 0.15   beta0 = 20.36   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.34562+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7}   kt2 = -0.02   at = 40500.0   ute = -1.613   ua1 = 1.0e-9   ub1 = -1.1724e-17   uc1 = -2.5133e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.745e-6   sbref = 1.74e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










* .model sky130_fd_pr__nfet_03v3_nvt__model.8 nmos  lmin = 5.95e-07 lmax = 6.05e-07 wmin = 6.95e-07 wmax = 7.05e-7   level = 54.0   tnom = 30.0   version = 4.5   toxm = 1.16e-8   xj = 1.5e-7   lln = 1.0   lwn = 1.0   wln = 1.0   wwn = 1.0   lint = {0+sky130_fd_pr__nfet_03v3_nvt__lint_diff}   ll = 0.0   lw = 0.0   lwl = 0.0   wint = {0+sky130_fd_pr__nfet_03v3_nvt__wint_diff}   wl = 0.0   ww = 0.0   wwl = 0.0   xl = 0.0   xw = 0.0   mobmod = 0.0   binunit = 2.0   dwg = 0.0   dwb = 0.0   igcmod = 0.0   igbmod = 0.0   rgatemod = 0.0   rbodymod = 1.0   trnqsmod = 0.0   acnqsmod = 0.0   fnoimod = 1.0   tnoimod = 1.0   permod = 1.0   geomod = 0.0   rdsmod = 0.0   tempmod = 0.0   lintnoi = 0.0   vfbsdoff = 0.0   lambda = 0.0   vtl = 0.0   lc = 5.0e-9   xn = 3.0   rnoia = 0.89   rnoib = 0.38   tnoia = 6.4e+6   tnoib = 7.2e+6   epsrox = 3.9   toxe = {1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.16e-008*sky130_fd_pr__nfet_03v3_nvt__toxe_mult*(sky130_fd_pr__nfet_03v3_nvt__toxe_slope/sqrt(l*w*mult)))}   dtox = 0.0   ndep = 1.7e+17   nsd = 1.0e+20   rshg = 0.1   rsh = {1*sky130_fd_pr__nfet_03v3_nvt__rshn_mult}   vth0 = {0.071092+sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__vth0_slope/sqrt(l*w*mult))}   k1 = 0.33502   k2 = {0+sky130_fd_pr__nfet_03v3_nvt__k2_diff_8}   k3 = 0.0   dvt0 = 1.0e-10   dvt1 = 0.536   dvt2 = -0.05   dvt0w = 0.0   dvt1w = 5000000.0   dvt2w = -0.032   w0 = 0.0   k3b = 0.0   phin = 0.01855708   lpe0 = -1.0e-10   lpeb = 0.0   vbm = -3.0   dvtp0 = 0.0   dvtp1 = 0.0   vsat = {120770+sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8}   ua = {4.145e-009+sky130_fd_pr__nfet_03v3_nvt__ua_diff_8}   ub = {3.7798e-019+sky130_fd_pr__nfet_03v3_nvt__ub_diff_8}   uc = 1.3541e-10   rdsw = {0+sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8}   prwb = 0.0   prwg = 0.0   wr = 1.0   u0 = {0.083529+sky130_fd_pr__nfet_03v3_nvt__u0_diff_8}   a0 = {0.00031139121+sky130_fd_pr__nfet_03v3_nvt__a0_diff_8}   keta = {0.0047834+sky130_fd_pr__nfet_03v3_nvt__keta_diff_8}   a1 = 0.0   a2 = 0.6218093   ags = {0.00014554757+sky130_fd_pr__nfet_03v3_nvt__ags_diff_8}   b0 = {0+sky130_fd_pr__nfet_03v3_nvt__b0_diff_8}   b1 = {0+sky130_fd_pr__nfet_03v3_nvt__b1_diff_8}   eu = 1.67   rdswmin = 0.0   rdw = 0.0   rdwmin = 0.0   rsw = 0.0   rswmin = 0.0   voff = {-0.098774+sky130_fd_pr__nfet_03v3_nvt__voff_diff_8+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__voff_slope/sqrt(l*w*mult))}   nfactor = {0.77345+sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_03v3_nvt__nfactor_slope/sqrt(l*w*mult))}   up = 0.0   ud = 0.0   lp = 1.0   tvfbsdoff = 0.0   tvoff = {0+sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8}   cit = -3.3686011e-37   cdsc = 0.0   cdscb = -0.0001   cdscd = 1.5e-5   eta0 = {0+sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8}   etab = 0.0   dsub = 0.071143   voffl = -2.9752837e-11   minv = 0.0   pclm = {2.8944111+sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8}   pdiblc1 = 0.87012255   pdiblc2 = 0.032974   pdiblcb = -0.05   drout = 0.27268   pscbe1 = 4.24e+9   pscbe2 = 1.0e-8   pvag = 5.2718232   delta = 0.01   alpha0 = 3.498e-7   alpha1 = 0.35   beta0 = 21.582   fprout = 10.125   pdits = {5.666761e-016+sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8}   pditsl = 0.0   pditsd = {0+sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8}   agidl = 0.0   bgidl = 2.3e+9   cgidl = 0.8   egidl = 0.5   aigbacc = 0.43   bigbacc = 0.054   cigbacc = 0.075   nigbacc = 1.0   aigbinv = 0.35   bigbinv = 0.03   cigbinv = 0.006   eigbinv = 1.1   nigbinv = 3.0   aigc = 0.43   bigc = 0.054   cigc = 0.075   nigc = 1.0   aigsd = 0.43   bigsd = 0.054   cigsd = 0.075   dlcig = 0.0   poxedge = 1.0   pigcd = 1.0   ntox = 1.0   toxref = 1.16e-8   kt1 = {-0.30496+sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8}   kt2 = -0.02   at = 34830.0   ute = -1.6817   ua1 = 1.0e-9   ub1 = -9.9403e-18   uc1 = -2.5133e-10   kt1l = 0.0   prt = 0.0   xrcrg1 = 12.0   xrcrg2 = 1.0   rbpb = 50.0   rbpd = 50.0   rbps = 50.0   rbdb = 50.0   rbsb = 50.0   gbmin = 1.0e-12   noia = 2.5e+41   noib = 0.0   noic = 0.0   em = 4.1000000e+7   af = 1.0   ef = 1.0   kf = 0.0   ntnoi = 1.0   dmcg = 0.0   dmcgt = 0.0   dmdg = 0.0   xgw = 0.0   xgl = 0.0   ngcon = 1.0   diomod = 1.0   njs = 1.5764   jss = 0.00042966   jsws = 8.040000000000001e-10   xtis = 0.0   bvs = 12.69   xjbvs = 1.0   ijthsrev = 0.1   ijthsfwd = 0.1   tpb = 0.0019685   tpbsw = 0.001   tpbswg = 0.0   tcj = 0.00083   tcjsw = 0.0   tcjswg = 0.0   cgdo = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgso = {3.2646e-010*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgbo = 0.0   capmod = 2.0   xpart = 0.0   cgsl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cgdl = {5e-011*sky130_fd_pr__nfet_03v3_nvt__overlap_mult}   cf = 0.0   clc = 1.0e-7   cle = 0.6   dlc = {6.5233e-008+sky130_fd_pr__nfet_03v3_nvt__dlc_diff+sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak}   dwc = {0+sky130_fd_pr__nfet_03v3_nvt__dwc_diff}   vfbcv = -1.0   acde = 0.4   moin = 15.0   noff = 4.00   voffcv = -0.14208   ngate = 1.0e+23   lwc = 0.0   llc = 0.0   lwlc = 0.0   wlc = 0.0   wwc = 0.0   wwlc = 0.0   ckappas = 0.6   cjs = {0.0008602*sky130_fd_pr__nfet_03v3_nvt__ajunction_mult}   mjs = 0.28329   pbs = 0.66345   cjsws = {8.5152e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjsws = 0.057926   pbsws = 1.0   cjswgs = {3.58e-011*sky130_fd_pr__nfet_03v3_nvt__pjunction_mult}   mjswgs = 0.33   pbswgs = 0.2442   saref = 1.95e-6   sbref = 1.94e-6   wlod = {0+sky130_fd_pr__nfet_03v3_nvt__wlod_diff}   kvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__kvth0_diff}   lkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff}   wkvth0 = {0+sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff}   pkvth0 = 0.0   llodvth = 0.0   wlodvth = 1.0   stk2 = 0.0   lodk2 = 1.0   lodeta0 = 1.0   ku0 = {0+sky130_fd_pr__nfet_03v3_nvt__ku0_diff}   lku0 = {0+sky130_fd_pr__nfet_03v3_nvt__lku0_diff}   wku0 = {0+sky130_fd_pr__nfet_03v3_nvt__wku0_diff}   pku0 = 0.0   llodku0 = 0.0   wlodku0 = 1.0   kvsat = {0+sky130_fd_pr__nfet_03v3_nvt__kvsat_diff}   steta0 = 0.0   tku0 = 0.0; HSpice Parser Retained (as a comment). Continuing.





















* DC IV MOS Parameters
* BSIM4 - Model Selectors
























* BSIM4 - Process Parameters






















* Threshold Voltage Parameters







* NEW BSIM4 Parameters for Level 54












* Mobility Parameters






* BSIM4 - Mobility Parameters
















* Subthreshold Current Parameters






* BSIM4 - Sub-threshold parameters














* Rout Parameters


* BSIM4 - Rout Parameters












* BSIM4 - Gate Induced Drain Leakage Model Parameters




* BSIM4 - Gate Leakage Current Parameters




* Temperature Effects Parameters





















* BSIM4 - High Speed RF Model Parameters









* BSIM4 - Flicker and Thermal Noise Parameters








* BSIM4 - Layout Dependent Parasitic Model Parameters








* Diode DC IV Parameters






* BSIM4 - Diode DC IV parameters
* Diode and FET Capacitance Parameters









* BSIM4 - FET and Diode capacitance parameters






























* Stress Parameters










.ENDS sky130_fd_pr__nfet_03v3_nvt





















