** Translated using xdm 2.6.0 on Nov_14_2022_16_05_28_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15 d g s b sky130_fd_pr__rf_nfet_01v8_bM02 w = 1.65 l = 0.15 m = 2 ad = 0.231 pd = 1.93 as = 0.462 ps = 3.86 nrd = 72.80 nrs = 36.40 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02 w = 1.65 l = 0.15 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 36.40 nrs = 0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15 d g s b sky130_fd_pr__rf_nfet_01v8_bM04 w = 1.65 l = 0.15 m = 4 ad = 0.231 pd = 1.93 as = 0.347 ps = 2.90 nrd = 72.80 nrs = 48.53 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04 w = 1.65 l = 0.15 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 36.40 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18 d g s b sky130_fd_pr__rf_nfet_01v8_bM02 w = 1.65 l = 0.18 m = 2 ad = 0.231 pd = 1.93 as = 0.462 ps = 3.86 nrd = 72.80 nrs = 36.40 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02 w = 1.65 l = 0.18 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 36.40 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18 d g s b sky130_fd_pr__rf_nfet_01v8_bM04 w = 1.65 l = 0.18 m = 4 ad = 0.231 pd = 1.93 as = 0.347 ps = 2.90 nrd = 72.80 nrs = 48.53 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04 w = 1.65 l = 0.18 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 36.40 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25 d g s b sky130_fd_pr__rf_nfet_01v8_bM02 w = 1.65 l = 0.25 m = 2 ad = 0.231 pd = 1.93 as = 0.462 ps = 3.86 nrd = 72.80 nrs = 36.40 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02 w = 1.65 l = 0.25 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 36.4 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25 d g s b sky130_fd_pr__rf_nfet_01v8_bM04 w = 1.65 l = 0.25 m = 4 ad = 0.231 pd = 1.93 as = 0.347 ps = 2.90 nrd = 72.80 nrs = 48.53 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04 w = 1.65 l = 0.25 m = 2 ad = 0.495 pd = 3.9 as = 0.0 ps = 0.0 nrd = 36.4 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15 d g s b sky130_fd_pr__rf_nfet_01v8_bM02W3p00 l = 0.15 m = 2 ad = 0.421 pd = 3.29 as = 0.843 ps = 6.58 nrd = 40.44 nrs = 20.22 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02W3p00 l = 0.15 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15 d g s b sky130_fd_pr__rf_nfet_01v8_bM04W3p00 l = 0.15 m = 4 ad = 0.421 pd = 3.29 as = 0.632 ps = 4.94 nrd = 40.44 nrs = 26.96 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04W3p00 l = 0.15 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18 d g s b sky130_fd_pr__rf_nfet_01v8_bM02W3p00 l = 0.18 m = 2 ad = 0.421 pd = 3.29 as = 0.843 ps = 6.58 nrd = 40.44 nrs = 20.22 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02W3p00 l = 0.18 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18 d g s b sky130_fd_pr__rf_nfet_01v8_bM04W3p00 l = 0.18 m = 4 ad = 0.421 pd = 3.29 as = 0.632 ps = 4.94 nrd = 40.44 nrs = 26.96 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04W3p00 l = 0.18 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25 d g s b sky130_fd_pr__rf_nfet_01v8_bM02W3p00 l = 0.25 m = 2 ad = 0.421 pd = 3.29 as = 0.843 ps = 6.58 nrd = 40.44 nrs = 20.22 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02W3p00 l = 0.25 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25 d g s b sky130_fd_pr__rf_nfet_01v8_bM04W3p00 l = 0.25 m = 4 ad = 0.421 pd = 3.29 as = 0.632 ps = 4.94 nrd = 40.44 nrs = 26.96 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04W3p00 l = 0.25 m = 2 ad = 0.903 pd = 6.62 as = 0.0 ps = 0.0 nrd = 20.22 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15 d g s b sky130_fd_pr__rf_nfet_01v8_bM02W5p00 l = 0.15 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 24.27 nrs = 12.13 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02W5p00 l = 0.15 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15 d g s b sky130_fd_pr__rf_nfet_01v8_bM04W5p00 l = 0.15 m = 4 ad = 0.707 pd = 5.33 as = 1.061 ps = 8.00 nrd = 24.27 nrs = 16.18 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04W5p00 l = 0.15 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18 d g s b sky130_fd_pr__rf_nfet_01v8_bM02W5p00 l = 0.18 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 24.27 nrs = 12.13 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02W5p00 l = 0.18 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18 d g s b sky130_fd_pr__rf_nfet_01v8_bM04W5p00 l = 0.18 m = 4 ad = 0.707 pd = 5.33 as = 1.061 ps = 8.00 nrd = 24.27 nrs = 16.18 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04W5p00 l = 0.18 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25 d g s b sky130_fd_pr__rf_nfet_01v8_bM02W5p00 l = 0.25 m = 2 ad = 0.707 pd = 5.33 as = 1.414 ps = 10.66 nrd = 24.27 nrs = 12.13 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM02W5p00 l = 0.25 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.0 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25
.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25 d g s b
.PARAM MULT=1.0

* xsky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25 d g s b sky130_fd_pr__rf_nfet_01v8_bM04W5p00 l = 0.25 m = 4 ad = 0.707 pd = 5.33 as = 1.061 ps = 8.00 nrd = 24.27 nrs = 16.18 mult = {4*mult}; HSpice Parser Retained (as a comment). Continuing.
* xsky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25_dummy b b s b sky130_fd_pr__rf_nfet_01v8_bM04W5p00 l = 0.25 m = 2 ad = 1.515 pd = 10.7 as = 0.0 ps = 0.00 nrd = 12.13 nrs = 0.0 mult = {2*mult}; HSpice Parser Retained (as a comment). Continuing.
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25
