** Translated using xdm 2.6.0 on Nov_14_2022_16_05_04_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE=3.689e-03
.PARAM SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE1=1.489e-02
.PARAM SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE2=1.689e-02
.PARAM SKY130_FD_PR__PFET_01V8_LVT__TOXE_SLOPE3=2.389e-02
.PARAM SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE=1.389e-02
.PARAM SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE1=9.789e-03
.PARAM SKY130_FD_PR__PFET_01V8_LVT__VTH0_SLOPE2=1.089e-02
.PARAM SKY130_FD_PR__PFET_01V8_LVT__LINT_SLOPE=0
.PARAM SKY130_FD_PR__PFET_01V8_LVT__WINT_SLOPE=0
.PARAM SKY130_FD_PR__PFET_01V8_LVT__NFACTOR_SLOPE=0.0
.PARAM SKY130_FD_PR__PFET_01V8_LVT__VOFF_SLOPE=0.0
