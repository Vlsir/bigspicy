** Translated using xdm 2.6.0 on Nov_14_2022_16_05_26_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

.PARAM SKY130_FD_PR__NPN_05V5_W1P00L2P00__IS_SLOPE_SPECTRE=0.0
.PARAM SKY130_FD_PR__NPN_05V5_W1P00L2P00__BF_SLOPE_SPECTRE=0.0
* statistics {
*   mismatch {
*     vary  sky130_fd_pr__npn_05v5_W1p00L2p00__is_slope_spectre dist=gauss std=1.0
*     vary  sky130_fd_pr__npn_05v5_W1p00L2p00__bf_slope_spectre dist=gauss std=1.0
*   }
* }
.SUBCKT sky130_fd_pr__npn_05v5_W1p00L2p00 c b e s
.PARAM MULT=1 AREA=1.0

Qsky130_fd_pr__npn_05v5_W1p00L2p00 c b e s 
+ sky130_fd_pr__npn_05v5_W1p00L2p00__model
* General Parameters
* Capacitance Parameters

* Noise Parameters





* DC Parameters

* Temperature Parameters






.ENDS sky130_fd_pr__npn_05v5_W1p00L2p00

















