** Translated using xdm 2.6.0 on Nov_14_2022_16_05_18_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 8
.PARAM 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TOXE_MULT=0.958 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RSHP_MULT=1.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__OVERLAP_MULT=0.7713 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AJUNCTION_MULT=9.5405e-1 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PJUNCTION_MULT=9.6374e-1 SKY130_FD_PR__ESD_PFET_G5V0D10V5__LINT_DIFF=1.21275e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__WINT_DIFF=-2.252e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__DLC_DIFF=1.21275e-8 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__DWC_DIFF=-2.252e-8 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_0=-0.001863 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_0=0.001058 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_0=-31427.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_0=0.041954 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_0=-0.08688 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_0=4.3035e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_0=-3.1175e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_0=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_0=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_0=0.021424 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_1=0.013438 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_1=-0.0020179 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_1=0.0010444 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_1=-28354.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_1=0.048874 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_1=-1.42e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_1=-0.065937 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_1=-2.3727e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_1=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_1=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_2=0.017194 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_2=-0.0016532 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_2=0.00075934 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_2=0.051024 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_2=-7.6179e-12 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_2=-27569.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_2=-0.094908 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_2=-2.0807e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_2=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_3=0.018257 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_3=-0.0025581 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_3=0.00124927 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_3=0.044703 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_3=7.5609e-12 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_3=-35289.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_3=-0.086391 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_3=-3.2769e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_3=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_4=0.025977 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_4=-0.0013669 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_4=0.00091382 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_4=0.043787 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_4=1.574e-10 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_4=-24808.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_4=0.078325 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_4=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_4=-4.9963e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_4=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_5=0.020181 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_5=-0.0021503 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_5=0.0010663 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_5=0.043391 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_5=-1.0798e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_5=-22995.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_5=-0.11963 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_5=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_5=-1.3111e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_6=-1.868e-19 SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_6=0.019337 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_6=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_6=-0.0018306 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_6=0.00086193 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_6=0.045188 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_6=-1.1042e-11 SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_6=-24982.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_6=-0.11297 SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_6=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__ETA0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UB_DIFF_7=-2.3793e-19 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__RDSW_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KETA_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__CGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__TVOFF_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__BGIDL_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITSD_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PCLM_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__AGIDL_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VOFF_DIFF_7=0.022032 SKY130_FD_PR__ESD_PFET_G5V0D10V5__A0_DIFF_7=0.0 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B0_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__K2_DIFF_7=-0.0019486 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__PDITS_DIFF_7=0.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__U0_DIFF_7=0.00096865 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VTH0_DIFF_7=0.045761 SKY130_FD_PR__ESD_PFET_G5V0D10V5__UA_DIFF_7=-2.12e-11 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__VSAT_DIFF_7=-21171.0 SKY130_FD_PR__ESD_PFET_G5V0D10V5__NFACTOR_DIFF_7=-0.13265 
+ SKY130_FD_PR__ESD_PFET_G5V0D10V5__B1_DIFF_7=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
*




* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
*























* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
.INCLUDE sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice























