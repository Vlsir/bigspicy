** Translated using xdm 2.6.0 on Nov_14_2022_16_05_20_PM
** from /tmp/_MEItbfi7Y/hspice.xml
** to /tmp/_MEItbfi7Y/xyce.xml

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SKY130 Spice File.

* Number of bins: 9
.PARAM 
+ SKY130_FD_PR__NFET_03V3_NVT__TOXE_MULT=0.9635 SKY130_FD_PR__NFET_03V3_NVT__RSHN_MULT=1.0 
+ SKY130_FD_PR__NFET_03V3_NVT__OVERLAP_MULT=0.51025 SKY130_FD_PR__NFET_03V3_NVT__AJUNCTION_MULT=0.68772 
+ SKY130_FD_PR__NFET_03V3_NVT__PJUNCTION_MULT=0.9019 SKY130_FD_PR__NFET_03V3_NVT__LINT_DIFF=1.21275e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__WINT_DIFF=-2.252e-8 SKY130_FD_PR__NFET_03V3_NVT__DLC_DIFF=1.6112e-8 
+ SKY130_FD_PR__NFET_03V3_NVT__DWC_DIFF=-2.252e-8 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_0=0.017139 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_0=-0.016856 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_0=-1.0949 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_0=-0.041263 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_0=0.00079908 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_0=-1877.8 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_0=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_0=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_0=-8.8355e-20 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_0=1.2237e-11 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_1=3.5287e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_1=0.010252 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_1=-0.00051272 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_1=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_1=-1.3847 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_1=-0.0485 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_1=-7.0468e-5 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_1=-9793.6 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_1=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_1=2.2579e-19 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_2=1.2013e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_2=1.1421e-10 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_2=0.0012159 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_2=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_2=-0.49031 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_2=-0.034235 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_2=0.0043842 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_2=-8139.1 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_2=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_3=6.5751e-20 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_3=2.2944e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_3=0.0177 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_3=-0.01428 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_3=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_3=-1.0283 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_3=-0.04376 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_3=0.0014903 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_3=-3761.4 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_3=0.0 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_4=-4.2142e-19 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_4=-1.3052e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_4=0.044934 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_4=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_4=0.0083971 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_4=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_4=-1.5502 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_4=-0.068861 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_4=0.0016304 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_4=-6110.3 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_5=0.01509 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_5=-5015.2 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_5=2.0257e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_5=4.4064e-11 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_5=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_5=0.0059498 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_5=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_5=-1.6314 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_5=0.014604 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_6=-0.77252 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_6=-0.0039098 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_6=0.011371 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_6=-3438.4 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_6=1.7785e-18 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_6=5.037e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_6=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_6=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_6=0.0058775 SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_7=0.021791 
+ SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_7=0.0022917 SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_7=-1.3041 SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_7=-0.046002 
+ SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_7=0.00087134 SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_7=-9538.4 
+ SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_7=4.1235e-19 
+ SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_7=2.4503e-11 
+ SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_7=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_7=0.0 SKY130_FD_PR__NFET_03V3_NVT__A0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PDITS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__TVOFF_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__VOFF_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__B0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__AGS_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__K2_DIFF_8=0.0038297 
+ SKY130_FD_PR__NFET_03V3_NVT__KT1_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__NFACTOR_DIFF_8=-0.51817 
+ SKY130_FD_PR__NFET_03V3_NVT__VTH0_DIFF_8=-0.040702 SKY130_FD_PR__NFET_03V3_NVT__U0_DIFF_8=0.006163 
+ SKY130_FD_PR__NFET_03V3_NVT__VSAT_DIFF_8=-7789.7 SKY130_FD_PR__NFET_03V3_NVT__B1_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UB_DIFF_8=1.381e-18 SKY130_FD_PR__NFET_03V3_NVT__ETA0_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__UA_DIFF_8=1.3573e-10 SKY130_FD_PR__NFET_03V3_NVT__KETA_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__RDSW_DIFF_8=0.0 SKY130_FD_PR__NFET_03V3_NVT__PDITSD_DIFF_8=0.0 
+ SKY130_FD_PR__NFET_03V3_NVT__PCLM_DIFF_8=0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
*














* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
*




















* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
.INCLUDE sky130_fd_pr__nfet_03v3_nvt.pm3.spice




















